module tt_um_rebeccargb_hardware_utf8 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_0_clk;
 wire retry;
 wire \u8.empty ;
 wire \u8.hs[0] ;
 wire \u8.hs[1] ;
 wire \u8.hs[2] ;
 wire \u8.hs[3] ;
 wire \u8.hs[4] ;
 wire \u8.hs[5] ;
 wire \u8.ls[0] ;
 wire \u8.ls[1] ;
 wire \u8.ls[2] ;
 wire \u8.ls[3] ;
 wire \u8.ls[4] ;
 wire \u8.ls[5] ;
 wire \u8.ls[6] ;
 wire \u8.ls[7] ;
 wire \u8.ls[8] ;
 wire \u8.ls[9] ;
 wire \u8.rbop[0] ;
 wire \u8.rbop[1] ;
 wire \u8.rbop[2] ;
 wire \u8.rc[16] ;
 wire \u8.rc[17] ;
 wire \u8.rc[18] ;
 wire \u8.rc[19] ;
 wire \u8.rc[20] ;
 wire \u8.rc[21] ;
 wire \u8.rc[22] ;
 wire \u8.rc[23] ;
 wire \u8.rc[24] ;
 wire \u8.rc[25] ;
 wire \u8.rc[26] ;
 wire \u8.rc[27] ;
 wire \u8.rc[28] ;
 wire \u8.rc[29] ;
 wire \u8.rc[30] ;
 wire \u8.rc[31] ;
 wire \u8.rcip[0] ;
 wire \u8.rcip[1] ;
 wire \u8.rcip[2] ;
 wire \u8.rcop[0] ;
 wire \u8.rcop[1] ;
 wire \u8.rcop[2] ;
 wire \u8.ruop[0] ;
 wire \u8.ruop[1] ;
 wire \u8.ruop[2] ;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;

 sg13g2_inv_1 _1073_ (.Y(_0188_),
    .A(net338));
 sg13g2_inv_4 _1074_ (.A(net341),
    .Y(_0189_));
 sg13g2_inv_4 _1075_ (.A(net342),
    .Y(_0190_));
 sg13g2_inv_4 _1076_ (.A(net343),
    .Y(_0191_));
 sg13g2_inv_1 _1077_ (.Y(_0192_),
    .A(net345));
 sg13g2_inv_4 _1078_ (.A(net346),
    .Y(_0193_));
 sg13g2_inv_4 _1079_ (.A(net348),
    .Y(_0194_));
 sg13g2_inv_1 _1080_ (.Y(_0195_),
    .A(\u8.ruop[2] ));
 sg13g2_inv_2 _1081_ (.Y(_0196_),
    .A(\u8.ruop[0] ));
 sg13g2_inv_2 _1082_ (.Y(_0197_),
    .A(net82));
 sg13g2_inv_1 _1083_ (.Y(_0198_),
    .A(\u8.rcip[0] ));
 sg13g2_inv_2 _1084_ (.Y(_0199_),
    .A(net349));
 sg13g2_inv_2 _1085_ (.Y(_0200_),
    .A(net355));
 sg13g2_inv_4 _1086_ (.A(net356),
    .Y(_0201_));
 sg13g2_inv_2 _1087_ (.Y(_0202_),
    .A(net357));
 sg13g2_inv_4 _1088_ (.A(net360),
    .Y(_0203_));
 sg13g2_inv_2 _1089_ (.Y(_0204_),
    .A(net369));
 sg13g2_inv_4 _1090_ (.A(net370),
    .Y(_0205_));
 sg13g2_inv_2 _1091_ (.Y(_0206_),
    .A(net371));
 sg13g2_inv_4 _1092_ (.A(\u8.ls[3] ),
    .Y(_0207_));
 sg13g2_inv_1 _1093_ (.Y(_0208_),
    .A(net373));
 sg13g2_inv_2 _1094_ (.Y(_0209_),
    .A(net374));
 sg13g2_inv_2 _1095_ (.Y(_0210_),
    .A(\u8.ls[0] ));
 sg13g2_inv_2 _1096_ (.Y(_0211_),
    .A(net375));
 sg13g2_inv_4 _1097_ (.A(net376),
    .Y(_0212_));
 sg13g2_inv_2 _1098_ (.Y(_0213_),
    .A(net378));
 sg13g2_inv_1 _1099_ (.Y(_0214_),
    .A(\u8.rc[28] ));
 sg13g2_inv_1 _1100_ (.Y(_0215_),
    .A(net106));
 sg13g2_inv_4 _1101_ (.A(net381),
    .Y(_0216_));
 sg13g2_inv_2 _1102_ (.Y(_0217_),
    .A(net382));
 sg13g2_inv_1 _1103_ (.Y(_0218_),
    .A(net7));
 sg13g2_inv_1 _1104_ (.Y(_0219_),
    .A(net14));
 sg13g2_inv_2 _1105_ (.Y(_0220_),
    .A(net15));
 sg13g2_inv_1 _1106_ (.Y(_0221_),
    .A(net10));
 sg13g2_inv_2 _1107_ (.Y(_0222_),
    .A(net400));
 sg13g2_inv_1 _1108_ (.Y(_0223_),
    .A(net11));
 sg13g2_inv_1 _1109_ (.Y(_0224_),
    .A(net12));
 sg13g2_inv_1 _1110_ (.Y(_0225_),
    .A(net2));
 sg13g2_inv_1 _1111_ (.Y(_0226_),
    .A(net8));
 sg13g2_inv_1 _1112_ (.Y(_0227_),
    .A(net9));
 sg13g2_nand2_1 _1113_ (.Y(_0228_),
    .A(net350),
    .B(net352));
 sg13g2_nor3_1 _1114_ (.A(_0201_),
    .B(_0202_),
    .C(_0228_),
    .Y(_0229_));
 sg13g2_nor3_1 _1115_ (.A(net338),
    .B(net339),
    .C(net340),
    .Y(_0230_));
 sg13g2_nor2_1 _1116_ (.A(net381),
    .B(net382),
    .Y(_0231_));
 sg13g2_or2_1 _1117_ (.X(_0232_),
    .B(net382),
    .A(\u8.rc[25] ));
 sg13g2_nor3_1 _1118_ (.A(\u8.rc[26] ),
    .B(net381),
    .C(net382),
    .Y(_0233_));
 sg13g2_and2_1 _1119_ (.A(_0230_),
    .B(_0233_),
    .X(_0234_));
 sg13g2_nor2_1 _1120_ (.A(\u8.rc[28] ),
    .B(net380),
    .Y(_0235_));
 sg13g2_and3_1 _1121_ (.X(_0236_),
    .A(_0230_),
    .B(_0233_),
    .C(_0235_));
 sg13g2_nand3_1 _1122_ (.B(_0233_),
    .C(_0235_),
    .A(_0230_),
    .Y(_0237_));
 sg13g2_nor2_1 _1123_ (.A(net346),
    .B(net347),
    .Y(_0238_));
 sg13g2_nor3_2 _1124_ (.A(net345),
    .B(net346),
    .C(net347),
    .Y(_0239_));
 sg13g2_nor4_1 _1125_ (.A(net342),
    .B(net343),
    .C(net378),
    .D(net379),
    .Y(_0240_));
 sg13g2_and3_2 _1126_ (.X(_0241_),
    .A(_0236_),
    .B(_0239_),
    .C(_0240_));
 sg13g2_nand3_1 _1127_ (.B(net351),
    .C(net354),
    .A(net349),
    .Y(_0242_));
 sg13g2_nand2_2 _1128_ (.Y(_0243_),
    .A(_0241_),
    .B(_0242_));
 sg13g2_nand2b_2 _1129_ (.Y(_0244_),
    .B(_0242_),
    .A_N(_0229_));
 sg13g2_nor3_1 _1130_ (.A(net377),
    .B(_0229_),
    .C(_0243_),
    .Y(_0245_));
 sg13g2_and2_1 _1131_ (.A(_0191_),
    .B(_0239_),
    .X(_0246_));
 sg13g2_or2_1 _1132_ (.X(_0247_),
    .B(\u8.rc[26] ),
    .A(net380));
 sg13g2_or4_1 _1133_ (.A(net376),
    .B(net378),
    .C(net379),
    .D(\u8.rc[28] ),
    .X(_0248_));
 sg13g2_nor4_1 _1134_ (.A(net376),
    .B(net378),
    .C(net379),
    .D(\u8.rc[26] ),
    .Y(_0249_));
 sg13g2_and4_1 _1135_ (.A(_0230_),
    .B(_0231_),
    .C(_0235_),
    .D(_0249_),
    .X(_0250_));
 sg13g2_or4_1 _1136_ (.A(net338),
    .B(net339),
    .C(net340),
    .D(net342),
    .X(_0251_));
 sg13g2_nor4_2 _1137_ (.A(_0232_),
    .B(_0247_),
    .C(_0248_),
    .Y(_0252_),
    .D(_0251_));
 sg13g2_and2_1 _1138_ (.A(_0246_),
    .B(_0252_),
    .X(_0253_));
 sg13g2_nand2_2 _1139_ (.Y(_0254_),
    .A(_0246_),
    .B(_0252_));
 sg13g2_nor2_2 _1140_ (.A(_0201_),
    .B(_0242_),
    .Y(_0255_));
 sg13g2_nand4_1 _1141_ (.B(net351),
    .C(net354),
    .A(net349),
    .Y(_0256_),
    .D(net356));
 sg13g2_nor2_1 _1142_ (.A(_0202_),
    .B(_0203_),
    .Y(_0257_));
 sg13g2_nand3_1 _1143_ (.B(net359),
    .C(net361),
    .A(net357),
    .Y(_0258_));
 sg13g2_nor2b_1 _1144_ (.A(net362),
    .B_N(net363),
    .Y(_0259_));
 sg13g2_and4_1 _1145_ (.A(net366),
    .B(net368),
    .C(_0257_),
    .D(_0259_),
    .X(_0260_));
 sg13g2_o21ai_1 _1146_ (.B1(_0260_),
    .Y(_0261_),
    .A1(net370),
    .A2(net371));
 sg13g2_a21oi_1 _1147_ (.A1(_0258_),
    .A2(_0261_),
    .Y(_0262_),
    .B1(_0256_));
 sg13g2_nand2b_1 _1148_ (.Y(_0263_),
    .B(_0253_),
    .A_N(_0262_));
 sg13g2_nor2_1 _1149_ (.A(_0205_),
    .B(_0206_),
    .Y(_0264_));
 sg13g2_nand2_1 _1150_ (.Y(_0265_),
    .A(net370),
    .B(net371));
 sg13g2_a22oi_1 _1151_ (.Y(_0266_),
    .B1(_0260_),
    .B2(_0264_),
    .A2(_0257_),
    .A1(net362));
 sg13g2_o21ai_1 _1152_ (.B1(_0253_),
    .Y(_0267_),
    .A1(_0256_),
    .A2(_0266_));
 sg13g2_nand4_1 _1153_ (.B(\u8.ls[3] ),
    .C(net373),
    .A(net368),
    .Y(_0268_),
    .D(net374));
 sg13g2_nor2_1 _1154_ (.A(_0265_),
    .B(_0268_),
    .Y(_0269_));
 sg13g2_nor2_1 _1155_ (.A(_0202_),
    .B(_0256_),
    .Y(_0270_));
 sg13g2_nand2_1 _1156_ (.Y(_0271_),
    .A(net357),
    .B(_0255_));
 sg13g2_nand2_1 _1157_ (.Y(_0272_),
    .A(net363),
    .B(net366));
 sg13g2_nand3_1 _1158_ (.B(net364),
    .C(net366),
    .A(net362),
    .Y(_0273_));
 sg13g2_nor3_2 _1159_ (.A(_0256_),
    .B(_0258_),
    .C(_0272_),
    .Y(_0274_));
 sg13g2_nand2_1 _1160_ (.Y(_0275_),
    .A(_0269_),
    .B(_0274_));
 sg13g2_nand2_1 _1161_ (.Y(_0276_),
    .A(net346),
    .B(net347));
 sg13g2_nand4_1 _1162_ (.B(net345),
    .C(net346),
    .A(net343),
    .Y(_0277_),
    .D(net347));
 sg13g2_nand4_1 _1163_ (.B(_0267_),
    .C(_0275_),
    .A(_0252_),
    .Y(_0278_),
    .D(_0277_));
 sg13g2_nand2_1 _1164_ (.Y(_0279_),
    .A(_0263_),
    .B(_0278_));
 sg13g2_nor2_1 _1165_ (.A(net361),
    .B(net364),
    .Y(_0280_));
 sg13g2_nor3_1 _1166_ (.A(net359),
    .B(net362),
    .C(net364),
    .Y(_0281_));
 sg13g2_o21ai_1 _1167_ (.B1(_0253_),
    .Y(_0282_),
    .A1(_0271_),
    .A2(_0281_));
 sg13g2_a21o_1 _1168_ (.A2(_0282_),
    .A1(_0279_),
    .B1(_0245_),
    .X(_0283_));
 sg13g2_nor4_1 _1169_ (.A(net351),
    .B(net354),
    .C(net356),
    .D(net357),
    .Y(_0284_));
 sg13g2_and2_1 _1170_ (.A(_0199_),
    .B(_0284_),
    .X(_0285_));
 sg13g2_nand4_1 _1171_ (.B(_0239_),
    .C(_0240_),
    .A(_0199_),
    .Y(_0286_),
    .D(_0284_));
 sg13g2_nor2_2 _1172_ (.A(_0237_),
    .B(_0286_),
    .Y(_0287_));
 sg13g2_nor4_1 _1173_ (.A(net359),
    .B(net362),
    .C(net363),
    .D(net365),
    .Y(_0288_));
 sg13g2_inv_1 _1174_ (.Y(_0289_),
    .A(_0288_));
 sg13g2_nor4_1 _1175_ (.A(net377),
    .B(_0237_),
    .C(_0286_),
    .D(_0289_),
    .Y(_0290_));
 sg13g2_nor3_1 _1176_ (.A(net366),
    .B(net368),
    .C(net370),
    .Y(_0291_));
 sg13g2_a21oi_1 _1177_ (.A1(\u8.ls[0] ),
    .A2(_0269_),
    .Y(_0292_),
    .B1(_0289_));
 sg13g2_nand3_1 _1178_ (.B(_0285_),
    .C(_0292_),
    .A(_0253_),
    .Y(_0293_));
 sg13g2_o21ai_1 _1179_ (.B1(net366),
    .Y(_0294_),
    .A1(net369),
    .A2(\u8.ls[5] ));
 sg13g2_a21o_1 _1180_ (.A2(_0294_),
    .A1(_0293_),
    .B1(_0291_),
    .X(_0295_));
 sg13g2_nand4_1 _1181_ (.B(_0281_),
    .C(_0287_),
    .A(_0212_),
    .Y(_0296_),
    .D(_0295_));
 sg13g2_nor3_2 _1182_ (.A(net375),
    .B(net377),
    .C(net2),
    .Y(_0297_));
 sg13g2_nand3_1 _1183_ (.B(_0296_),
    .C(_0297_),
    .A(_0283_),
    .Y(_0298_));
 sg13g2_nand3_1 _1184_ (.B(net378),
    .C(net379),
    .A(net376),
    .Y(_0299_));
 sg13g2_nand3_1 _1185_ (.B(net380),
    .C(\u8.rc[26] ),
    .A(\u8.rc[28] ),
    .Y(_0300_));
 sg13g2_nor4_2 _1186_ (.A(_0212_),
    .B(_0213_),
    .C(net379),
    .Y(_0301_),
    .D(_0300_));
 sg13g2_nor2_1 _1187_ (.A(_0190_),
    .B(_0191_),
    .Y(_0302_));
 sg13g2_a21oi_1 _1188_ (.A1(net342),
    .A2(net344),
    .Y(_0303_),
    .B1(net341));
 sg13g2_nand3_1 _1189_ (.B(net339),
    .C(net382),
    .A(net338),
    .Y(_0304_));
 sg13g2_o21ai_1 _1190_ (.B1(_0216_),
    .Y(_0305_),
    .A1(_0303_),
    .A2(_0304_));
 sg13g2_nand2_1 _1191_ (.Y(_0306_),
    .A(_0301_),
    .B(_0305_));
 sg13g2_nand2_1 _1192_ (.Y(_0307_),
    .A(_0299_),
    .B(_0306_));
 sg13g2_nor3_1 _1193_ (.A(_0299_),
    .B(_0300_),
    .C(_0304_),
    .Y(_0308_));
 sg13g2_nor4_2 _1194_ (.A(_0216_),
    .B(_0299_),
    .C(_0300_),
    .Y(_0309_),
    .D(_0304_));
 sg13g2_nand3_1 _1195_ (.B(net343),
    .C(net345),
    .A(net342),
    .Y(_0310_));
 sg13g2_nor3_1 _1196_ (.A(_0189_),
    .B(_0193_),
    .C(_0310_),
    .Y(_0311_));
 sg13g2_and2_1 _1197_ (.A(_0309_),
    .B(_0311_),
    .X(_0312_));
 sg13g2_nor3_1 _1198_ (.A(_0265_),
    .B(_0268_),
    .C(_0272_),
    .Y(_0313_));
 sg13g2_nand2b_1 _1199_ (.Y(_0314_),
    .B(net369),
    .A_N(_0313_));
 sg13g2_nor3_1 _1200_ (.A(_0189_),
    .B(_0276_),
    .C(_0310_),
    .Y(_0315_));
 sg13g2_and2_1 _1201_ (.A(_0309_),
    .B(_0315_),
    .X(_0316_));
 sg13g2_nand3_1 _1202_ (.B(net350),
    .C(net352),
    .A(net348),
    .Y(_0317_));
 sg13g2_and3_1 _1203_ (.X(_0318_),
    .A(_0274_),
    .B(_0309_),
    .C(_0315_));
 sg13g2_a21oi_1 _1204_ (.A1(_0314_),
    .A2(_0318_),
    .Y(_0319_),
    .B1(_0271_));
 sg13g2_or4_1 _1205_ (.A(_0189_),
    .B(_0299_),
    .C(_0300_),
    .D(_0304_),
    .X(_0320_));
 sg13g2_or4_1 _1206_ (.A(_0193_),
    .B(_0216_),
    .C(_0310_),
    .D(_0320_),
    .X(_0321_));
 sg13g2_or3_1 _1207_ (.A(_0194_),
    .B(_0242_),
    .C(_0321_),
    .X(_0322_));
 sg13g2_o21ai_1 _1208_ (.B1(_0316_),
    .Y(_0323_),
    .A1(_0319_),
    .A2(_0322_));
 sg13g2_nand2_1 _1209_ (.Y(_0324_),
    .A(_0302_),
    .B(_0323_));
 sg13g2_nand2_1 _1210_ (.Y(_0325_),
    .A(net340),
    .B(_0308_));
 sg13g2_a21oi_1 _1211_ (.A1(_0302_),
    .A2(_0323_),
    .Y(_0326_),
    .B1(_0325_));
 sg13g2_a21oi_1 _1212_ (.A1(_0189_),
    .A2(_0310_),
    .Y(_0327_),
    .B1(_0304_));
 sg13g2_o21ai_1 _1213_ (.B1(_0301_),
    .Y(_0328_),
    .A1(net381),
    .A2(_0327_));
 sg13g2_nor4_1 _1214_ (.A(_0194_),
    .B(net355),
    .C(_0203_),
    .D(\u8.rc[25] ),
    .Y(_0329_));
 sg13g2_nor3_1 _1215_ (.A(net341),
    .B(net346),
    .C(_0280_),
    .Y(_0330_));
 sg13g2_and4_1 _1216_ (.A(_0244_),
    .B(_0301_),
    .C(_0329_),
    .D(_0330_),
    .X(_0331_));
 sg13g2_nor3_1 _1217_ (.A(_0201_),
    .B(_0258_),
    .C(_0317_),
    .Y(_0332_));
 sg13g2_nor2b_1 _1218_ (.A(_0332_),
    .B_N(_0327_),
    .Y(_0333_));
 sg13g2_a22oi_1 _1219_ (.Y(_0334_),
    .B1(_0331_),
    .B2(_0333_),
    .A2(_0328_),
    .A1(_0299_));
 sg13g2_nor3_1 _1220_ (.A(\u8.rc[25] ),
    .B(_0299_),
    .C(_0300_),
    .Y(_0335_));
 sg13g2_nand2b_1 _1221_ (.Y(_0336_),
    .B(_0334_),
    .A_N(_0335_));
 sg13g2_o21ai_1 _1222_ (.B1(_0307_),
    .Y(_0337_),
    .A1(_0326_),
    .A2(_0336_));
 sg13g2_nor2_1 _1223_ (.A(net375),
    .B(_0225_),
    .Y(_0338_));
 sg13g2_nand2_1 _1224_ (.Y(_0339_),
    .A(net337),
    .B(_0337_));
 sg13g2_o21ai_1 _1225_ (.B1(_0298_),
    .Y(uo_out[0]),
    .A1(_0225_),
    .A2(_0339_));
 sg13g2_nor2b_1 _1226_ (.A(_0296_),
    .B_N(_0297_),
    .Y(_0340_));
 sg13g2_a21o_2 _1227_ (.A2(net2),
    .A1(retry),
    .B1(_0340_),
    .X(uo_out[1]));
 sg13g2_and4_1 _1228_ (.A(net376),
    .B(net378),
    .C(net379),
    .D(\u8.rc[28] ),
    .X(_0341_));
 sg13g2_nand4_1 _1229_ (.B(net378),
    .C(net379),
    .A(net376),
    .Y(_0342_),
    .D(\u8.rc[28] ));
 sg13g2_nand2_1 _1230_ (.Y(_0343_),
    .A(net380),
    .B(_0341_));
 sg13g2_and4_1 _1231_ (.A(_0189_),
    .B(_0190_),
    .C(_0191_),
    .D(_0239_),
    .X(_0344_));
 sg13g2_nand2_1 _1232_ (.Y(_0345_),
    .A(_0194_),
    .B(_0285_));
 sg13g2_nand4_1 _1233_ (.B(_0255_),
    .C(_0288_),
    .A(_0202_),
    .Y(_0346_),
    .D(_0316_));
 sg13g2_nand2_1 _1234_ (.Y(_0347_),
    .A(_0345_),
    .B(_0346_));
 sg13g2_a21o_1 _1235_ (.A2(_0347_),
    .A1(_0312_),
    .B1(_0344_),
    .X(_0348_));
 sg13g2_or2_1 _1236_ (.X(_0349_),
    .B(_0348_),
    .A(_0324_));
 sg13g2_o21ai_1 _1237_ (.B1(_0308_),
    .Y(_0350_),
    .A1(net340),
    .A2(_0344_));
 sg13g2_nand2b_1 _1238_ (.Y(_0351_),
    .B(_0349_),
    .A_N(_0350_));
 sg13g2_nor2_1 _1239_ (.A(_0234_),
    .B(_0335_),
    .Y(_0352_));
 sg13g2_a21oi_1 _1240_ (.A1(_0351_),
    .A2(_0352_),
    .Y(_0353_),
    .B1(_0343_));
 sg13g2_o21ai_1 _1241_ (.B1(_0334_),
    .Y(_0354_),
    .A1(_0247_),
    .A2(_0342_));
 sg13g2_o21ai_1 _1242_ (.B1(_0307_),
    .Y(_0355_),
    .A1(_0353_),
    .A2(_0354_));
 sg13g2_nand3_1 _1243_ (.B(_0338_),
    .C(_0355_),
    .A(net377),
    .Y(_0356_));
 sg13g2_o21ai_1 _1244_ (.B1(_0297_),
    .Y(_0357_),
    .A1(_0229_),
    .A2(_0243_));
 sg13g2_o21ai_1 _1245_ (.B1(_0356_),
    .Y(uo_out[2]),
    .A1(_0243_),
    .A2(_0357_));
 sg13g2_a21oi_1 _1246_ (.A1(_0309_),
    .A2(_0348_),
    .Y(_0358_),
    .B1(_0234_));
 sg13g2_o21ai_1 _1247_ (.B1(_0247_),
    .Y(_0359_),
    .A1(_0343_),
    .A2(_0358_));
 sg13g2_nand3_1 _1248_ (.B(_0341_),
    .C(_0359_),
    .A(_0338_),
    .Y(_0360_));
 sg13g2_nand2_1 _1249_ (.Y(_0361_),
    .A(_0200_),
    .B(_0203_));
 sg13g2_a21oi_2 _1250_ (.B1(_0254_),
    .Y(_0362_),
    .A2(_0361_),
    .A1(_0244_));
 sg13g2_o21ai_1 _1251_ (.B1(_0250_),
    .Y(_0363_),
    .A1(_0190_),
    .A2(_0246_));
 sg13g2_and2_1 _1252_ (.A(net3),
    .B(_0363_),
    .X(_0364_));
 sg13g2_nor2_1 _1253_ (.A(_0253_),
    .B(_0364_),
    .Y(_0365_));
 sg13g2_nor2_1 _1254_ (.A(_0362_),
    .B(_0365_),
    .Y(_0366_));
 sg13g2_o21ai_1 _1255_ (.B1(_0360_),
    .Y(uo_out[3]),
    .A1(_0357_),
    .A2(_0366_));
 sg13g2_nor3_1 _1256_ (.A(net375),
    .B(net377),
    .C(_0225_),
    .Y(_0367_));
 sg13g2_nand2_1 _1257_ (.Y(_0368_),
    .A(_0363_),
    .B(_0367_));
 sg13g2_a22oi_1 _1258_ (.Y(_0369_),
    .B1(_0277_),
    .B2(_0252_),
    .A2(_0274_),
    .A1(_0269_));
 sg13g2_nand2b_1 _1259_ (.Y(_0370_),
    .B(_0369_),
    .A_N(_0364_));
 sg13g2_nand2_1 _1260_ (.Y(_0371_),
    .A(_0282_),
    .B(_0370_));
 sg13g2_a21oi_1 _1261_ (.A1(_0243_),
    .A2(_0371_),
    .Y(_0372_),
    .B1(_0362_));
 sg13g2_a21oi_1 _1262_ (.A1(net353),
    .A2(net355),
    .Y(_0373_),
    .B1(net359));
 sg13g2_nand3_1 _1263_ (.B(_0273_),
    .C(_0373_),
    .A(_0241_),
    .Y(_0374_));
 sg13g2_nand2b_1 _1264_ (.Y(_0375_),
    .B(_0374_),
    .A_N(_0357_));
 sg13g2_o21ai_1 _1265_ (.B1(_0368_),
    .Y(uo_out[4]),
    .A1(_0372_),
    .A2(_0375_));
 sg13g2_o21ai_1 _1266_ (.B1(_0267_),
    .Y(_0376_),
    .A1(_0275_),
    .A2(_0364_));
 sg13g2_nand3_1 _1267_ (.B(_0297_),
    .C(_0376_),
    .A(_0263_),
    .Y(_0377_));
 sg13g2_a22oi_1 _1268_ (.Y(_0378_),
    .B1(_0364_),
    .B2(_0367_),
    .A2(net2),
    .A1(retry));
 sg13g2_nand4_1 _1269_ (.B(_0360_),
    .C(_0377_),
    .A(_0356_),
    .Y(uo_out[5]),
    .D(_0378_));
 sg13g2_nor3_2 _1270_ (.A(\u8.empty ),
    .B(_0253_),
    .C(_0363_),
    .Y(_0379_));
 sg13g2_nand3b_1 _1271_ (.B(_0254_),
    .C(_0211_),
    .Y(_0380_),
    .A_N(_0363_));
 sg13g2_nand4_1 _1272_ (.B(_0301_),
    .C(_0305_),
    .A(_0299_),
    .Y(_0381_),
    .D(_0328_));
 sg13g2_nand2_1 _1273_ (.Y(_0382_),
    .A(_0254_),
    .B(_0381_));
 sg13g2_a21oi_2 _1274_ (.B1(net375),
    .Y(_0383_),
    .A2(_0381_),
    .A1(_0254_));
 sg13g2_a21o_1 _1275_ (.A2(_0381_),
    .A1(_0254_),
    .B1(net375),
    .X(_0384_));
 sg13g2_nor2_1 _1276_ (.A(\u8.ruop[1] ),
    .B(net313),
    .Y(_0385_));
 sg13g2_nand2_1 _1277_ (.Y(_0386_),
    .A(net337),
    .B(_0307_));
 sg13g2_nor2_2 _1278_ (.A(_0334_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_a21o_1 _1279_ (.A2(_0387_),
    .A1(_0196_),
    .B1(_0385_),
    .X(_0388_));
 sg13g2_a22oi_1 _1280_ (.Y(_0389_),
    .B1(net313),
    .B2(\u8.ruop[1] ),
    .A2(_0380_),
    .A1(\u8.ruop[2] ));
 sg13g2_a22oi_1 _1281_ (.Y(_0390_),
    .B1(_0388_),
    .B2(_0389_),
    .A2(net320),
    .A1(_0195_));
 sg13g2_nand2_1 _1282_ (.Y(_0391_),
    .A(net399),
    .B(net301));
 sg13g2_o21ai_1 _1283_ (.B1(_0391_),
    .Y(uo_out[6]),
    .A1(net399),
    .A2(_0380_));
 sg13g2_a22oi_1 _1284_ (.Y(_0392_),
    .B1(_0309_),
    .B2(_0311_),
    .A2(_0252_),
    .A1(_0246_));
 sg13g2_nand2_1 _1285_ (.Y(_0393_),
    .A(net376),
    .B(_0342_));
 sg13g2_a21oi_1 _1286_ (.A1(net376),
    .A2(_0342_),
    .Y(_0394_),
    .B1(net375));
 sg13g2_nand2_1 _1287_ (.Y(_0395_),
    .A(net337),
    .B(_0393_));
 sg13g2_nand2_2 _1288_ (.Y(_0396_),
    .A(_0392_),
    .B(net335));
 sg13g2_or2_1 _1289_ (.X(_0397_),
    .B(_0318_),
    .A(_0290_));
 sg13g2_a22oi_1 _1290_ (.Y(_0398_),
    .B1(_0341_),
    .B2(net380),
    .A2(_0249_),
    .A1(_0235_));
 sg13g2_nand2_1 _1291_ (.Y(_0399_),
    .A(_0393_),
    .B(_0398_));
 sg13g2_and2_1 _1292_ (.A(_0392_),
    .B(_0399_),
    .X(_0400_));
 sg13g2_a221oi_1 _1293_ (.B2(_0399_),
    .C1(_0290_),
    .B1(_0392_),
    .A1(_0274_),
    .Y(_0401_),
    .A2(_0316_));
 sg13g2_nand2_1 _1294_ (.Y(_0402_),
    .A(net337),
    .B(_0401_));
 sg13g2_or3_1 _1295_ (.A(_0236_),
    .B(_0309_),
    .C(_0398_),
    .X(_0403_));
 sg13g2_a221oi_1 _1296_ (.B2(_0403_),
    .C1(_0287_),
    .B1(_0392_),
    .A1(_0255_),
    .Y(_0404_),
    .A2(_0316_));
 sg13g2_nor4_2 _1297_ (.A(net375),
    .B(_0397_),
    .C(_0400_),
    .Y(_0405_),
    .D(_0404_));
 sg13g2_nand2b_2 _1298_ (.Y(_0406_),
    .B(_0405_),
    .A_N(net319));
 sg13g2_nand2b_1 _1299_ (.Y(_0407_),
    .B(_0406_),
    .A_N(net398));
 sg13g2_and2_1 _1300_ (.A(\u8.rbop[2] ),
    .B(net319),
    .X(_0408_));
 sg13g2_or2_1 _1301_ (.X(_0409_),
    .B(net319),
    .A(\u8.rbop[2] ));
 sg13g2_nor2_1 _1302_ (.A(\u8.rbop[1] ),
    .B(_0402_),
    .Y(_0410_));
 sg13g2_xor2_1 _1303_ (.B(_0402_),
    .A(\u8.rbop[1] ),
    .X(_0411_));
 sg13g2_o21ai_1 _1304_ (.B1(net337),
    .Y(_0412_),
    .A1(_0397_),
    .A2(_0404_));
 sg13g2_nand2_1 _1305_ (.Y(_0413_),
    .A(\u8.rbop[0] ),
    .B(net312));
 sg13g2_a21oi_1 _1306_ (.A1(_0411_),
    .A2(_0413_),
    .Y(_0414_),
    .B1(_0410_));
 sg13g2_o21ai_1 _1307_ (.B1(_0409_),
    .Y(_0415_),
    .A1(_0408_),
    .A2(_0414_));
 sg13g2_nor2_1 _1308_ (.A(\u8.rbop[0] ),
    .B(net312),
    .Y(_0416_));
 sg13g2_xor2_1 _1309_ (.B(net312),
    .A(\u8.rbop[0] ),
    .X(_0417_));
 sg13g2_nand2_1 _1310_ (.Y(_0418_),
    .A(_0411_),
    .B(_0417_));
 sg13g2_nand3_1 _1311_ (.B(_0411_),
    .C(_0417_),
    .A(_0409_),
    .Y(_0419_));
 sg13g2_nand3_1 _1312_ (.B(net300),
    .C(_0419_),
    .A(net398),
    .Y(_0420_));
 sg13g2_and2_1 _1313_ (.A(_0407_),
    .B(_0420_),
    .X(uo_out[7]));
 sg13g2_or2_1 _1314_ (.X(_0421_),
    .B(net312),
    .A(_0401_));
 sg13g2_nor2_2 _1315_ (.A(net319),
    .B(_0421_),
    .Y(_0422_));
 sg13g2_or3_1 _1316_ (.A(net319),
    .B(_0401_),
    .C(net312),
    .X(_0423_));
 sg13g2_a21oi_2 _1317_ (.B1(net319),
    .Y(_0424_),
    .A2(_0401_),
    .A1(net337));
 sg13g2_nand2_1 _1318_ (.Y(_0425_),
    .A(\u8.rc[18] ),
    .B(net311));
 sg13g2_and3_2 _1319_ (.X(_0426_),
    .A(net337),
    .B(_0401_),
    .C(_0404_));
 sg13g2_and2_1 _1320_ (.A(net319),
    .B(_0405_),
    .X(_0427_));
 sg13g2_and2_1 _1321_ (.A(net312),
    .B(net311),
    .X(_0428_));
 sg13g2_a221oi_1 _1322_ (.B2(net311),
    .C1(_0426_),
    .B1(net312),
    .A1(net319),
    .Y(_0429_),
    .A2(_0405_));
 sg13g2_and2_1 _1323_ (.A(_0423_),
    .B(_0429_),
    .X(_0430_));
 sg13g2_a21oi_1 _1324_ (.A1(_0280_),
    .A2(_0291_),
    .Y(_0431_),
    .B1(net359));
 sg13g2_and4_1 _1325_ (.A(net347),
    .B(_0270_),
    .C(_0312_),
    .D(_0431_),
    .X(_0432_));
 sg13g2_inv_2 _1326_ (.Y(_0433_),
    .A(_0432_));
 sg13g2_and4_1 _1327_ (.A(net346),
    .B(_0396_),
    .C(_0405_),
    .D(_0433_),
    .X(_0434_));
 sg13g2_a21oi_1 _1328_ (.A1(_0203_),
    .A2(_0284_),
    .Y(_0435_),
    .B1(net349));
 sg13g2_nand2_1 _1329_ (.Y(_0436_),
    .A(_0316_),
    .B(_0435_));
 sg13g2_nand3_1 _1330_ (.B(_0426_),
    .C(_0436_),
    .A(net343),
    .Y(_0437_));
 sg13g2_nand2b_2 _1331_ (.Y(_0438_),
    .B(_0437_),
    .A_N(_0434_));
 sg13g2_nor2_2 _1332_ (.A(net307),
    .B(_0438_),
    .Y(_0439_));
 sg13g2_nor4_1 _1333_ (.A(net371),
    .B(\u8.ls[3] ),
    .C(net373),
    .D(net374),
    .Y(_0440_));
 sg13g2_nor3_1 _1334_ (.A(_0204_),
    .B(\u8.ls[5] ),
    .C(_0440_),
    .Y(_0441_));
 sg13g2_nand4_1 _1335_ (.B(_0274_),
    .C(_0312_),
    .A(net348),
    .Y(_0442_),
    .D(_0441_));
 sg13g2_nand2_1 _1336_ (.Y(_0443_),
    .A(\u8.rc[18] ),
    .B(net316));
 sg13g2_a22oi_1 _1337_ (.Y(_0444_),
    .B1(_0443_),
    .B2(net308),
    .A2(_0439_),
    .A1(_0425_));
 sg13g2_nor2_2 _1338_ (.A(net399),
    .B(net7),
    .Y(_0445_));
 sg13g2_nand2_1 _1339_ (.Y(_0446_),
    .A(net395),
    .B(_0445_));
 sg13g2_nand3_1 _1340_ (.B(net334),
    .C(_0445_),
    .A(net395),
    .Y(_0447_));
 sg13g2_inv_1 _1341_ (.Y(_0448_),
    .A(_0447_));
 sg13g2_nor2_2 _1342_ (.A(net399),
    .B(net395),
    .Y(_0449_));
 sg13g2_or2_1 _1343_ (.X(_0450_),
    .B(net395),
    .A(net399));
 sg13g2_a21o_2 _1344_ (.A2(net324),
    .A1(_0220_),
    .B1(_0446_),
    .X(_0451_));
 sg13g2_a21oi_2 _1345_ (.B1(_0446_),
    .Y(_0452_),
    .A2(net324),
    .A1(_0220_));
 sg13g2_o21ai_1 _1346_ (.B1(net315),
    .Y(_0453_),
    .A1(net325),
    .A2(_0444_));
 sg13g2_nand2_1 _1347_ (.Y(_0454_),
    .A(_0219_),
    .B(net15));
 sg13g2_nand2b_1 _1348_ (.Y(_0455_),
    .B(_0339_),
    .A_N(_0454_));
 sg13g2_a221oi_1 _1349_ (.B2(_0429_),
    .C1(_0454_),
    .B1(_0421_),
    .A1(net337),
    .Y(_0456_),
    .A2(_0337_));
 sg13g2_nor2_1 _1350_ (.A(_0447_),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_nor2_1 _1351_ (.A(_0445_),
    .B(net387),
    .Y(_0458_));
 sg13g2_a21oi_2 _1352_ (.B1(net399),
    .Y(_0459_),
    .A2(net7),
    .A1(net5));
 sg13g2_nor2_1 _1353_ (.A(net399),
    .B(net6),
    .Y(_0460_));
 sg13g2_o21ai_1 _1354_ (.B1(net1),
    .Y(_0461_),
    .A1(_0459_),
    .A2(_0460_));
 sg13g2_a21oi_1 _1355_ (.A1(\u8.rcip[2] ),
    .A2(net390),
    .Y(_0462_),
    .B1(_0461_));
 sg13g2_nand2_1 _1356_ (.Y(_0463_),
    .A(_0458_),
    .B(_0460_));
 sg13g2_nor2_1 _1357_ (.A(net313),
    .B(_0387_),
    .Y(_0464_));
 sg13g2_nand2b_1 _1358_ (.Y(_0465_),
    .B(_0383_),
    .A_N(_0387_));
 sg13g2_o21ai_1 _1359_ (.B1(_0462_),
    .Y(_0466_),
    .A1(_0380_),
    .A2(_0463_));
 sg13g2_a21oi_1 _1360_ (.A1(_0244_),
    .A2(_0362_),
    .Y(_0467_),
    .B1(_0463_));
 sg13g2_a21oi_1 _1361_ (.A1(net306),
    .A2(_0467_),
    .Y(_0468_),
    .B1(_0466_));
 sg13g2_nor2b_2 _1362_ (.A(_0457_),
    .B_N(_0468_),
    .Y(_0469_));
 sg13g2_o21ai_1 _1363_ (.B1(_0468_),
    .Y(_0470_),
    .A1(_0447_),
    .A2(_0456_));
 sg13g2_nor2_2 _1364_ (.A(\u8.rcip[2] ),
    .B(_0450_),
    .Y(_0471_));
 sg13g2_nand2_2 _1365_ (.Y(_0472_),
    .A(net82),
    .B(_0471_));
 sg13g2_nor2_2 _1366_ (.A(_0198_),
    .B(_0472_),
    .Y(_0473_));
 sg13g2_nor2_2 _1367_ (.A(net348),
    .B(net393),
    .Y(_0474_));
 sg13g2_o21ai_1 _1368_ (.B1(net323),
    .Y(_0475_),
    .A1(net409),
    .A2(net8));
 sg13g2_nor2_2 _1369_ (.A(net320),
    .B(_0383_),
    .Y(_0476_));
 sg13g2_nand2_2 _1370_ (.Y(_0477_),
    .A(_0380_),
    .B(net313));
 sg13g2_nor2_2 _1371_ (.A(_0387_),
    .B(_0477_),
    .Y(_0478_));
 sg13g2_o21ai_1 _1372_ (.B1(_0458_),
    .Y(_0479_),
    .A1(net305),
    .A2(_0478_));
 sg13g2_o21ai_1 _1373_ (.B1(_0479_),
    .Y(_0480_),
    .A1(_0474_),
    .A2(_0475_));
 sg13g2_nor2_1 _1374_ (.A(_0470_),
    .B(_0480_),
    .Y(_0481_));
 sg13g2_o21ai_1 _1375_ (.B1(net416),
    .Y(_0482_),
    .A1(net98),
    .A2(_0469_));
 sg13g2_a21oi_1 _1376_ (.A1(_0453_),
    .A2(_0481_),
    .Y(_0000_),
    .B1(_0482_));
 sg13g2_nand2_1 _1377_ (.Y(_0483_),
    .A(net344),
    .B(net316));
 sg13g2_nand2_1 _1378_ (.Y(_0484_),
    .A(net344),
    .B(net311));
 sg13g2_a22oi_1 _1379_ (.Y(_0485_),
    .B1(_0484_),
    .B2(_0439_),
    .A2(_0483_),
    .A1(net307));
 sg13g2_o21ai_1 _1380_ (.B1(net315),
    .Y(_0486_),
    .A1(net325),
    .A2(_0485_));
 sg13g2_nand2_1 _1381_ (.Y(_0487_),
    .A(_0193_),
    .B(net409));
 sg13g2_nor2_1 _1382_ (.A(net412),
    .B(net9),
    .Y(_0488_));
 sg13g2_nand2_1 _1383_ (.Y(_0489_),
    .A(net393),
    .B(_0227_));
 sg13g2_nand3_1 _1384_ (.B(_0487_),
    .C(_0489_),
    .A(net323),
    .Y(_0490_));
 sg13g2_nand2_1 _1385_ (.Y(_0491_),
    .A(_0486_),
    .B(_0490_));
 sg13g2_o21ai_1 _1386_ (.B1(net416),
    .Y(_0492_),
    .A1(_0470_),
    .A2(_0491_));
 sg13g2_a21oi_1 _1387_ (.A1(_0216_),
    .A2(_0470_),
    .Y(_0001_),
    .B1(_0492_));
 sg13g2_nand2_1 _1388_ (.Y(_0493_),
    .A(net342),
    .B(net311));
 sg13g2_nand2_1 _1389_ (.Y(_0494_),
    .A(\u8.rc[20] ),
    .B(net316));
 sg13g2_a22oi_1 _1390_ (.Y(_0495_),
    .B1(_0494_),
    .B2(net307),
    .A2(_0493_),
    .A1(_0439_));
 sg13g2_o21ai_1 _1391_ (.B1(_0452_),
    .Y(_0496_),
    .A1(net324),
    .A2(_0495_));
 sg13g2_nor2_2 _1392_ (.A(\u8.rc[18] ),
    .B(net394),
    .Y(_0497_));
 sg13g2_nor2_1 _1393_ (.A(net10),
    .B(net412),
    .Y(_0498_));
 sg13g2_or4_1 _1394_ (.A(_0198_),
    .B(_0472_),
    .C(_0497_),
    .D(_0498_),
    .X(_0499_));
 sg13g2_nand3_1 _1395_ (.B(_0496_),
    .C(_0499_),
    .A(_0479_),
    .Y(_0500_));
 sg13g2_o21ai_1 _1396_ (.B1(net417),
    .Y(_0501_),
    .A1(_0470_),
    .A2(_0500_));
 sg13g2_a21oi_1 _1397_ (.A1(_0215_),
    .A2(_0470_),
    .Y(_0002_),
    .B1(_0501_));
 sg13g2_a21oi_1 _1398_ (.A1(net307),
    .A2(net318),
    .Y(_0502_),
    .B1(_0422_));
 sg13g2_nand2_1 _1399_ (.Y(_0503_),
    .A(_0199_),
    .B(_0246_));
 sg13g2_nor2_1 _1400_ (.A(\u8.rc[20] ),
    .B(_0216_),
    .Y(_0504_));
 sg13g2_nand4_1 _1401_ (.B(_0308_),
    .C(_0503_),
    .A(net340),
    .Y(_0505_),
    .D(_0504_));
 sg13g2_and2_1 _1402_ (.A(_0428_),
    .B(_0505_),
    .X(_0506_));
 sg13g2_nand2_1 _1403_ (.Y(_0507_),
    .A(_0428_),
    .B(_0505_));
 sg13g2_a21oi_1 _1404_ (.A1(_0502_),
    .A2(_0507_),
    .Y(_0508_),
    .B1(_0189_));
 sg13g2_nor3_1 _1405_ (.A(net325),
    .B(_0438_),
    .C(_0508_),
    .Y(_0509_));
 sg13g2_or2_1 _1406_ (.X(_0510_),
    .B(_0509_),
    .A(_0451_));
 sg13g2_nand2_1 _1407_ (.Y(_0511_),
    .A(_0191_),
    .B(net403));
 sg13g2_nor2_1 _1408_ (.A(net412),
    .B(net11),
    .Y(_0512_));
 sg13g2_nand3b_1 _1409_ (.B(net323),
    .C(_0511_),
    .Y(_0513_),
    .A_N(_0512_));
 sg13g2_nand4_1 _1410_ (.B(_0479_),
    .C(_0510_),
    .A(net291),
    .Y(_0514_),
    .D(_0513_));
 sg13g2_o21ai_1 _1411_ (.B1(net416),
    .Y(_0515_),
    .A1(net380),
    .A2(net291));
 sg13g2_nor2b_1 _1412_ (.A(_0515_),
    .B_N(_0514_),
    .Y(_0003_));
 sg13g2_nand2_1 _1413_ (.Y(_0516_),
    .A(net339),
    .B(net318));
 sg13g2_o21ai_1 _1414_ (.B1(_0335_),
    .Y(_0517_),
    .A1(\u8.rc[24] ),
    .A2(_0251_));
 sg13g2_a221oi_1 _1415_ (.B2(_0422_),
    .C1(_0438_),
    .B1(_0517_),
    .A1(\u8.rc[24] ),
    .Y(_0518_),
    .A2(_0506_));
 sg13g2_nand2b_1 _1416_ (.Y(_0519_),
    .B(_0518_),
    .A_N(net307));
 sg13g2_a21oi_1 _1417_ (.A1(net339),
    .A2(_0422_),
    .Y(_0520_),
    .B1(_0519_));
 sg13g2_a21oi_1 _1418_ (.A1(net307),
    .A2(_0516_),
    .Y(_0521_),
    .B1(_0520_));
 sg13g2_o21ai_1 _1419_ (.B1(net315),
    .Y(_0522_),
    .A1(net325),
    .A2(_0521_));
 sg13g2_nor2_1 _1420_ (.A(_0190_),
    .B(net394),
    .Y(_0523_));
 sg13g2_nor2_1 _1421_ (.A(net409),
    .B(_0224_),
    .Y(_0524_));
 sg13g2_o21ai_1 _1422_ (.B1(_0473_),
    .Y(_0525_),
    .A1(_0523_),
    .A2(_0524_));
 sg13g2_and3_1 _1423_ (.X(_0526_),
    .A(net291),
    .B(_0479_),
    .C(_0525_));
 sg13g2_o21ai_1 _1424_ (.B1(net416),
    .Y(_0527_),
    .A1(net105),
    .A2(net291));
 sg13g2_a21oi_1 _1425_ (.A1(_0522_),
    .A2(_0526_),
    .Y(_0004_),
    .B1(_0527_));
 sg13g2_nand2_1 _1426_ (.Y(_0528_),
    .A(net338),
    .B(net318));
 sg13g2_and2_1 _1427_ (.A(net307),
    .B(_0528_),
    .X(_0529_));
 sg13g2_a21oi_1 _1428_ (.A1(net338),
    .A2(_0422_),
    .Y(_0530_),
    .B1(_0519_));
 sg13g2_o21ai_1 _1429_ (.B1(net335),
    .Y(_0531_),
    .A1(_0529_),
    .A2(_0530_));
 sg13g2_nor2_1 _1430_ (.A(net407),
    .B(net13),
    .Y(_0532_));
 sg13g2_a21oi_1 _1431_ (.A1(_0189_),
    .A2(net408),
    .Y(_0533_),
    .B1(_0532_));
 sg13g2_a22oi_1 _1432_ (.Y(_0534_),
    .B1(_0533_),
    .B2(net323),
    .A2(_0531_),
    .A1(net315));
 sg13g2_o21ai_1 _1433_ (.B1(net416),
    .Y(_0535_),
    .A1(net379),
    .A2(net291));
 sg13g2_a21oi_1 _1434_ (.A1(net291),
    .A2(_0534_),
    .Y(_0005_),
    .B1(_0535_));
 sg13g2_and2_1 _1435_ (.A(net335),
    .B(_0518_),
    .X(_0536_));
 sg13g2_o21ai_1 _1436_ (.B1(_0536_),
    .Y(_0537_),
    .A1(_0217_),
    .A2(_0502_));
 sg13g2_nor2_1 _1437_ (.A(net339),
    .B(net392),
    .Y(_0538_));
 sg13g2_nor2_1 _1438_ (.A(net14),
    .B(net407),
    .Y(_0539_));
 sg13g2_nor2_1 _1439_ (.A(_0538_),
    .B(_0539_),
    .Y(_0540_));
 sg13g2_a22oi_1 _1440_ (.Y(_0541_),
    .B1(_0540_),
    .B2(net323),
    .A2(_0537_),
    .A1(net315));
 sg13g2_nand3_1 _1441_ (.B(_0479_),
    .C(_0541_),
    .A(_0469_),
    .Y(_0542_));
 sg13g2_o21ai_1 _1442_ (.B1(net416),
    .Y(_0543_),
    .A1(net96),
    .A2(net291));
 sg13g2_nor2b_1 _1443_ (.A(_0543_),
    .B_N(_0542_),
    .Y(_0006_));
 sg13g2_nand2_1 _1444_ (.Y(_0544_),
    .A(_0212_),
    .B(_0470_));
 sg13g2_nand3_1 _1445_ (.B(net308),
    .C(net318),
    .A(net381),
    .Y(_0545_));
 sg13g2_nand2_1 _1446_ (.Y(_0546_),
    .A(_0536_),
    .B(_0545_));
 sg13g2_nor2_1 _1447_ (.A(_0220_),
    .B(net414),
    .Y(_0547_));
 sg13g2_a21o_1 _1448_ (.A2(net407),
    .A1(\u8.rc[23] ),
    .B1(_0547_),
    .X(_0548_));
 sg13g2_a22oi_1 _1449_ (.Y(_0549_),
    .B1(_0548_),
    .B2(net323),
    .A2(_0546_),
    .A1(net315));
 sg13g2_nand3_1 _1450_ (.B(_0479_),
    .C(_0549_),
    .A(net291),
    .Y(_0550_));
 sg13g2_and3_1 _1451_ (.X(_0007_),
    .A(net416),
    .B(_0544_),
    .C(_0550_));
 sg13g2_nor2_1 _1452_ (.A(net334),
    .B(_0446_),
    .Y(_0551_));
 sg13g2_and2_1 _1453_ (.A(net365),
    .B(net401),
    .X(_0552_));
 sg13g2_nand2b_1 _1454_ (.Y(_0553_),
    .B(net400),
    .A_N(net365));
 sg13g2_or2_1 _1455_ (.X(_0554_),
    .B(_0552_),
    .A(_0547_));
 sg13g2_nand2_1 _1456_ (.Y(_0555_),
    .A(_0205_),
    .B(net408));
 sg13g2_nand2b_2 _1457_ (.Y(_0556_),
    .B(_0555_),
    .A_N(_0532_));
 sg13g2_nand2_1 _1458_ (.Y(_0557_),
    .A(net372),
    .B(net411));
 sg13g2_nand2_1 _1459_ (.Y(_0558_),
    .A(_0206_),
    .B(net405));
 sg13g2_nor2b_2 _1460_ (.A(_0524_),
    .B_N(_0557_),
    .Y(_0559_));
 sg13g2_inv_1 _1461_ (.Y(_0560_),
    .A(_0559_));
 sg13g2_nor2_1 _1462_ (.A(net373),
    .B(net392),
    .Y(_0561_));
 sg13g2_nand2_2 _1463_ (.Y(_0562_),
    .A(_0208_),
    .B(net400));
 sg13g2_nand2b_2 _1464_ (.Y(_0563_),
    .B(_0562_),
    .A_N(_0498_));
 sg13g2_inv_1 _1465_ (.Y(_0564_),
    .A(_0563_));
 sg13g2_nand2_1 _1466_ (.Y(_0565_),
    .A(_0204_),
    .B(net405));
 sg13g2_a21oi_2 _1467_ (.B1(_0539_),
    .Y(_0566_),
    .A2(net407),
    .A1(_0204_));
 sg13g2_nand2_1 _1468_ (.Y(_0567_),
    .A(_0207_),
    .B(net402));
 sg13g2_a21oi_1 _1469_ (.A1(_0207_),
    .A2(net412),
    .Y(_0568_),
    .B1(_0512_));
 sg13g2_inv_1 _1470_ (.Y(_0569_),
    .A(_0568_));
 sg13g2_nand4_1 _1471_ (.B(_0556_),
    .C(_0566_),
    .A(_0554_),
    .Y(_0570_),
    .D(_0568_));
 sg13g2_nor3_2 _1472_ (.A(_0559_),
    .B(_0563_),
    .C(_0570_),
    .Y(_0571_));
 sg13g2_inv_2 _1473_ (.Y(_0572_),
    .A(_0571_));
 sg13g2_nand2_2 _1474_ (.Y(_0573_),
    .A(_0382_),
    .B(_0387_));
 sg13g2_inv_1 _1475_ (.Y(_0574_),
    .A(net302));
 sg13g2_nor2_2 _1476_ (.A(_0572_),
    .B(net302),
    .Y(_0575_));
 sg13g2_nand3_1 _1477_ (.B(_0387_),
    .C(_0571_),
    .A(_0382_),
    .Y(_0576_));
 sg13g2_nor4_1 _1478_ (.A(net4),
    .B(net6),
    .C(_0478_),
    .D(_0575_),
    .Y(_0577_));
 sg13g2_and3_1 _1479_ (.X(_0578_),
    .A(_0244_),
    .B(_0362_),
    .C(_0383_));
 sg13g2_o21ai_1 _1480_ (.B1(net302),
    .Y(_0579_),
    .A1(_0387_),
    .A2(_0578_));
 sg13g2_a21oi_1 _1481_ (.A1(_0577_),
    .A2(_0579_),
    .Y(_0580_),
    .B1(_0459_));
 sg13g2_o21ai_1 _1482_ (.B1(net1),
    .Y(_0581_),
    .A1(_0447_),
    .A2(_0455_));
 sg13g2_nor4_1 _1483_ (.A(_0471_),
    .B(_0551_),
    .C(_0580_),
    .D(_0581_),
    .Y(_0582_));
 sg13g2_o21ai_1 _1484_ (.B1(net416),
    .Y(_0583_),
    .A1(net97),
    .A2(_0582_));
 sg13g2_inv_1 _1485_ (.Y(_0008_),
    .A(_0583_));
 sg13g2_nor2b_2 _1486_ (.A(net395),
    .B_N(net396),
    .Y(_0584_));
 sg13g2_nand2b_2 _1487_ (.Y(_0585_),
    .B(net396),
    .A_N(net395));
 sg13g2_or2_1 _1488_ (.X(_0586_),
    .B(_0414_),
    .A(_0409_));
 sg13g2_nor2_1 _1489_ (.A(_0411_),
    .B(_0416_),
    .Y(_0587_));
 sg13g2_a21oi_2 _1490_ (.B1(_0587_),
    .Y(_0588_),
    .A2(_0413_),
    .A1(_0411_));
 sg13g2_and3_2 _1491_ (.X(_0589_),
    .A(net300),
    .B(net297),
    .C(_0588_));
 sg13g2_nor2b_2 _1492_ (.A(_0411_),
    .B_N(_0417_),
    .Y(_0590_));
 sg13g2_and3_2 _1493_ (.X(_0591_),
    .A(net300),
    .B(net297),
    .C(_0590_));
 sg13g2_nor3_2 _1494_ (.A(_0409_),
    .B(_0414_),
    .C(_0417_),
    .Y(_0592_));
 sg13g2_nor2_2 _1495_ (.A(_0409_),
    .B(_0418_),
    .Y(_0593_));
 sg13g2_or2_1 _1496_ (.X(_0594_),
    .B(_0593_),
    .A(_0592_));
 sg13g2_nor4_1 _1497_ (.A(_0210_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0595_));
 sg13g2_nand4_1 _1498_ (.B(net299),
    .C(net297),
    .A(net368),
    .Y(_0596_),
    .D(_0590_));
 sg13g2_nand4_1 _1499_ (.B(net299),
    .C(net297),
    .A(net356),
    .Y(_0597_),
    .D(_0588_));
 sg13g2_nor3_2 _1500_ (.A(\u8.rbop[2] ),
    .B(\u8.rbop[1] ),
    .C(\u8.rbop[0] ),
    .Y(_0598_));
 sg13g2_inv_2 _1501_ (.Y(_0599_),
    .A(_0598_));
 sg13g2_a22oi_1 _1502_ (.Y(_0600_),
    .B1(_0593_),
    .B2(net345),
    .A2(_0592_),
    .A1(net382));
 sg13g2_nand4_1 _1503_ (.B(_0597_),
    .C(_0599_),
    .A(_0596_),
    .Y(_0601_),
    .D(_0600_));
 sg13g2_nor2_1 _1504_ (.A(net7),
    .B(_0420_),
    .Y(_0602_));
 sg13g2_nand4_1 _1505_ (.B(_0218_),
    .C(net300),
    .A(net398),
    .Y(_0603_),
    .D(_0419_));
 sg13g2_and3_2 _1506_ (.X(_0604_),
    .A(_0406_),
    .B(_0423_),
    .C(_0429_));
 sg13g2_nand2_1 _1507_ (.Y(_0605_),
    .A(_0406_),
    .B(net308));
 sg13g2_nand2_1 _1508_ (.Y(_0606_),
    .A(_0212_),
    .B(net378));
 sg13g2_nand3_1 _1509_ (.B(_0412_),
    .C(net311),
    .A(net345),
    .Y(_0607_));
 sg13g2_o21ai_1 _1510_ (.B1(_0607_),
    .Y(_0608_),
    .A1(_0406_),
    .A2(_0606_));
 sg13g2_a221oi_1 _1511_ (.B2(net368),
    .C1(_0608_),
    .B1(_0427_),
    .A1(net382),
    .Y(_0609_),
    .A2(_0422_));
 sg13g2_a221oi_1 _1512_ (.B2(\u8.ls[0] ),
    .C1(_0599_),
    .B1(_0604_),
    .A1(net356),
    .Y(_0610_),
    .A2(_0426_));
 sg13g2_a21oi_1 _1513_ (.A1(_0609_),
    .A2(_0610_),
    .Y(_0611_),
    .B1(_0603_));
 sg13g2_o21ai_1 _1514_ (.B1(_0611_),
    .Y(_0612_),
    .A1(_0595_),
    .A2(_0601_));
 sg13g2_nor2_2 _1515_ (.A(net363),
    .B(net402),
    .Y(_0613_));
 sg13g2_nor2_1 _1516_ (.A(_0474_),
    .B(_0613_),
    .Y(_0614_));
 sg13g2_nor3_2 _1517_ (.A(\u8.ruop[2] ),
    .B(\u8.ruop[1] ),
    .C(_0196_),
    .Y(_0615_));
 sg13g2_or3_1 _1518_ (.A(\u8.ruop[2] ),
    .B(\u8.ruop[1] ),
    .C(_0196_),
    .X(_0616_));
 sg13g2_nor2b_2 _1519_ (.A(\u8.ruop[2] ),
    .B_N(\u8.ruop[1] ),
    .Y(_0617_));
 sg13g2_and2_1 _1520_ (.A(_0196_),
    .B(_0617_),
    .X(_0618_));
 sg13g2_or2_1 _1521_ (.X(_0619_),
    .B(net327),
    .A(net330));
 sg13g2_nor3_1 _1522_ (.A(_0474_),
    .B(_0613_),
    .C(_0619_),
    .Y(_0620_));
 sg13g2_nor2_1 _1523_ (.A(_0194_),
    .B(net403),
    .Y(_0621_));
 sg13g2_a21o_1 _1524_ (.A2(net403),
    .A1(net363),
    .B1(_0621_),
    .X(_0622_));
 sg13g2_a221oi_1 _1525_ (.B2(net331),
    .C1(_0620_),
    .B1(_0622_),
    .A1(\u8.ls[0] ),
    .Y(_0623_),
    .A2(net328));
 sg13g2_xnor2_1 _1526_ (.Y(_0624_),
    .A(net345),
    .B(_0238_));
 sg13g2_nor2_2 _1527_ (.A(net360),
    .B(net393),
    .Y(_0625_));
 sg13g2_a21oi_1 _1528_ (.A1(net391),
    .A2(_0624_),
    .Y(_0626_),
    .B1(_0625_));
 sg13g2_nand2_1 _1529_ (.Y(_0627_),
    .A(net331),
    .B(_0626_));
 sg13g2_nor2_2 _1530_ (.A(_0210_),
    .B(net409),
    .Y(_0628_));
 sg13g2_a21oi_1 _1531_ (.A1(net363),
    .A2(net404),
    .Y(_0629_),
    .B1(_0628_));
 sg13g2_nor2b_1 _1532_ (.A(_0629_),
    .B_N(net328),
    .Y(_0630_));
 sg13g2_nor2_2 _1533_ (.A(\u8.ls[0] ),
    .B(net393),
    .Y(_0631_));
 sg13g2_and2_1 _1534_ (.A(\u8.ruop[0] ),
    .B(_0617_),
    .X(_0632_));
 sg13g2_nand2_1 _1535_ (.Y(_0633_),
    .A(\u8.ruop[0] ),
    .B(_0617_));
 sg13g2_nor3_1 _1536_ (.A(_0613_),
    .B(_0631_),
    .C(_0633_),
    .Y(_0634_));
 sg13g2_nor2_2 _1537_ (.A(net332),
    .B(_0617_),
    .Y(_0635_));
 sg13g2_or2_1 _1538_ (.X(_0636_),
    .B(_0617_),
    .A(net332));
 sg13g2_nor3_1 _1539_ (.A(_0630_),
    .B(_0634_),
    .C(net322),
    .Y(_0637_));
 sg13g2_nor2_1 _1540_ (.A(net359),
    .B(net406),
    .Y(_0638_));
 sg13g2_a21o_1 _1541_ (.A2(_0624_),
    .A1(net402),
    .B1(_0638_),
    .X(_0639_));
 sg13g2_a22oi_1 _1542_ (.Y(_0640_),
    .B1(_0639_),
    .B2(net322),
    .A2(_0637_),
    .A1(_0627_));
 sg13g2_a21oi_1 _1543_ (.A1(net320),
    .A2(_0640_),
    .Y(_0641_),
    .B1(_0476_));
 sg13g2_o21ai_1 _1544_ (.B1(_0641_),
    .Y(_0642_),
    .A1(net302),
    .A2(_0623_));
 sg13g2_o21ai_1 _1545_ (.B1(net332),
    .Y(_0643_),
    .A1(_0613_),
    .A2(_0631_));
 sg13g2_a21oi_1 _1546_ (.A1(net329),
    .A2(_0629_),
    .Y(_0644_),
    .B1(net303));
 sg13g2_a21oi_1 _1547_ (.A1(_0643_),
    .A2(_0644_),
    .Y(_0645_),
    .B1(_0642_));
 sg13g2_nor2b_1 _1548_ (.A(net7),
    .B_N(net396),
    .Y(_0646_));
 sg13g2_nand2_2 _1549_ (.Y(_0647_),
    .A(net398),
    .B(_0218_));
 sg13g2_o21ai_1 _1550_ (.B1(_0647_),
    .Y(_0648_),
    .A1(\u8.ls[0] ),
    .A2(net309));
 sg13g2_or3_1 _1551_ (.A(net301),
    .B(_0645_),
    .C(_0648_),
    .X(_0649_));
 sg13g2_a21o_1 _1552_ (.A2(_0649_),
    .A1(_0612_),
    .B1(net385),
    .X(_0650_));
 sg13g2_nand2b_1 _1553_ (.Y(_0651_),
    .B(net396),
    .A_N(net6));
 sg13g2_and3_2 _1554_ (.X(_0652_),
    .A(_0585_),
    .B(_0647_),
    .C(_0651_));
 sg13g2_nand3_1 _1555_ (.B(_0647_),
    .C(_0651_),
    .A(_0585_),
    .Y(_0653_));
 sg13g2_nand2b_1 _1556_ (.Y(_0654_),
    .B(\u8.rcop[1] ),
    .A_N(\u8.rcop[2] ));
 sg13g2_nor2b_1 _1557_ (.A(net74),
    .B_N(net70),
    .Y(_0655_));
 sg13g2_nand2b_2 _1558_ (.Y(_0656_),
    .B(\u8.rcop[0] ),
    .A_N(\u8.rcop[2] ));
 sg13g2_and2_1 _1559_ (.A(\u8.rcop[1] ),
    .B(_0655_),
    .X(_0657_));
 sg13g2_nand2_1 _1560_ (.Y(_0658_),
    .A(net85),
    .B(_0655_));
 sg13g2_a21oi_1 _1561_ (.A1(_0217_),
    .A2(net394),
    .Y(_0659_),
    .B1(_0631_));
 sg13g2_and2_1 _1562_ (.A(_0654_),
    .B(_0656_),
    .X(_0660_));
 sg13g2_nor2_2 _1563_ (.A(\u8.rcop[1] ),
    .B(_0656_),
    .Y(_0661_));
 sg13g2_a22oi_1 _1564_ (.Y(_0662_),
    .B1(_0661_),
    .B2(_0614_),
    .A2(_0659_),
    .A1(_0657_));
 sg13g2_nor2_2 _1565_ (.A(\u8.rcop[0] ),
    .B(_0654_),
    .Y(_0663_));
 sg13g2_a21oi_1 _1566_ (.A1(_0622_),
    .A2(_0663_),
    .Y(_0664_),
    .B1(net326));
 sg13g2_nor2_2 _1567_ (.A(net74),
    .B(_0585_),
    .Y(_0665_));
 sg13g2_a21oi_1 _1568_ (.A1(net382),
    .A2(net403),
    .Y(_0666_),
    .B1(_0628_));
 sg13g2_a22oi_1 _1569_ (.Y(_0667_),
    .B1(_0666_),
    .B2(net326),
    .A2(_0664_),
    .A1(_0662_));
 sg13g2_a21oi_1 _1570_ (.A1(net336),
    .A2(_0667_),
    .Y(_0668_),
    .B1(_0652_));
 sg13g2_and2_1 _1571_ (.A(net1),
    .B(net421),
    .X(_0669_));
 sg13g2_nand2_2 _1572_ (.Y(_0670_),
    .A(net1),
    .B(net421));
 sg13g2_o21ai_1 _1573_ (.B1(net383),
    .Y(_0671_),
    .A1(net88),
    .A2(_0653_));
 sg13g2_a21oi_1 _1574_ (.A1(_0650_),
    .A2(_0668_),
    .Y(_0009_),
    .B1(_0671_));
 sg13g2_nor4_1 _1575_ (.A(_0209_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0672_));
 sg13g2_nand4_1 _1576_ (.B(net299),
    .C(net298),
    .A(net365),
    .Y(_0673_),
    .D(_0590_));
 sg13g2_nand4_1 _1577_ (.B(net299),
    .C(net298),
    .A(net354),
    .Y(_0674_),
    .D(_0588_));
 sg13g2_a22oi_1 _1578_ (.Y(_0675_),
    .B1(_0593_),
    .B2(net343),
    .A2(_0592_),
    .A1(net381));
 sg13g2_nand4_1 _1579_ (.B(_0673_),
    .C(_0674_),
    .A(_0599_),
    .Y(_0676_),
    .D(_0675_));
 sg13g2_nand2_1 _1580_ (.Y(_0677_),
    .A(net374),
    .B(_0604_));
 sg13g2_nand2_1 _1581_ (.Y(_0678_),
    .A(net365),
    .B(_0427_));
 sg13g2_a21oi_1 _1582_ (.A1(net354),
    .A2(_0426_),
    .Y(_0679_),
    .B1(_0599_));
 sg13g2_nand2_1 _1583_ (.Y(_0680_),
    .A(_0678_),
    .B(_0679_));
 sg13g2_a221oi_1 _1584_ (.B2(net343),
    .C1(_0680_),
    .B1(_0428_),
    .A1(net381),
    .Y(_0681_),
    .A2(_0422_));
 sg13g2_a21oi_1 _1585_ (.A1(_0677_),
    .A2(_0681_),
    .Y(_0682_),
    .B1(_0603_));
 sg13g2_o21ai_1 _1586_ (.B1(_0682_),
    .Y(_0683_),
    .A1(_0672_),
    .A2(_0676_));
 sg13g2_nor2_1 _1587_ (.A(net301),
    .B(_0646_),
    .Y(_0684_));
 sg13g2_o21ai_1 _1588_ (.B1(_0487_),
    .Y(_0685_),
    .A1(net361),
    .A2(net409));
 sg13g2_nor2_1 _1589_ (.A(net361),
    .B(net393),
    .Y(_0686_));
 sg13g2_a21oi_1 _1590_ (.A1(_0193_),
    .A2(net394),
    .Y(_0687_),
    .B1(_0686_));
 sg13g2_a22oi_1 _1591_ (.Y(_0688_),
    .B1(_0687_),
    .B2(net331),
    .A2(net328),
    .A1(net374));
 sg13g2_o21ai_1 _1592_ (.B1(_0688_),
    .Y(_0689_),
    .A1(_0619_),
    .A2(_0685_));
 sg13g2_xnor2_1 _1593_ (.Y(_0690_),
    .A(net343),
    .B(_0239_));
 sg13g2_nor2_2 _1594_ (.A(net358),
    .B(net393),
    .Y(_0691_));
 sg13g2_a21oi_1 _1595_ (.A1(net392),
    .A2(_0690_),
    .Y(_0692_),
    .B1(_0691_));
 sg13g2_nor2_1 _1596_ (.A(\u8.ls[1] ),
    .B(net410),
    .Y(_0693_));
 sg13g2_nor2_1 _1597_ (.A(_0686_),
    .B(_0693_),
    .Y(_0694_));
 sg13g2_nand2_2 _1598_ (.Y(_0695_),
    .A(_0209_),
    .B(net407));
 sg13g2_o21ai_1 _1599_ (.B1(_0695_),
    .Y(_0696_),
    .A1(net362),
    .A2(net403));
 sg13g2_o21ai_1 _1600_ (.B1(_0636_),
    .Y(_0697_),
    .A1(_0633_),
    .A2(_0696_));
 sg13g2_a221oi_1 _1601_ (.B2(net328),
    .C1(_0697_),
    .B1(_0694_),
    .A1(net332),
    .Y(_0698_),
    .A2(_0692_));
 sg13g2_nor2_1 _1602_ (.A(net357),
    .B(net402),
    .Y(_0699_));
 sg13g2_a21oi_1 _1603_ (.A1(net402),
    .A2(_0690_),
    .Y(_0700_),
    .B1(_0699_));
 sg13g2_o21ai_1 _1604_ (.B1(_0379_),
    .Y(_0701_),
    .A1(_0636_),
    .A2(_0700_));
 sg13g2_o21ai_1 _1605_ (.B1(net309),
    .Y(_0702_),
    .A1(_0698_),
    .A2(_0701_));
 sg13g2_nor2_1 _1606_ (.A(net332),
    .B(_0694_),
    .Y(_0703_));
 sg13g2_a21oi_1 _1607_ (.A1(net332),
    .A2(_0696_),
    .Y(_0704_),
    .B1(_0703_));
 sg13g2_a221oi_1 _1608_ (.B2(net306),
    .C1(_0702_),
    .B1(_0704_),
    .A1(_0574_),
    .Y(_0705_),
    .A2(_0689_));
 sg13g2_nor2_1 _1609_ (.A(net374),
    .B(net309),
    .Y(_0706_));
 sg13g2_or4_1 _1610_ (.A(net301),
    .B(_0646_),
    .C(_0705_),
    .D(_0706_),
    .X(_0707_));
 sg13g2_a21o_1 _1611_ (.A2(_0707_),
    .A1(_0683_),
    .B1(net385),
    .X(_0708_));
 sg13g2_nor3_1 _1612_ (.A(\u8.rcop[1] ),
    .B(_0656_),
    .C(_0685_),
    .Y(_0709_));
 sg13g2_a21oi_1 _1613_ (.A1(_0663_),
    .A2(_0687_),
    .Y(_0710_),
    .B1(_0709_));
 sg13g2_a21oi_1 _1614_ (.A1(_0216_),
    .A2(net404),
    .Y(_0711_),
    .B1(_0693_));
 sg13g2_o21ai_1 _1615_ (.B1(_0695_),
    .Y(_0712_),
    .A1(net381),
    .A2(net400));
 sg13g2_o21ai_1 _1616_ (.B1(_0710_),
    .Y(_0713_),
    .A1(_0658_),
    .A2(_0712_));
 sg13g2_a21oi_1 _1617_ (.A1(_0660_),
    .A2(_0711_),
    .Y(_0714_),
    .B1(_0713_));
 sg13g2_nor2b_1 _1618_ (.A(_0714_),
    .B_N(net336),
    .Y(_0715_));
 sg13g2_nor2_1 _1619_ (.A(_0652_),
    .B(_0715_),
    .Y(_0716_));
 sg13g2_o21ai_1 _1620_ (.B1(net384),
    .Y(_0717_),
    .A1(net87),
    .A2(_0653_));
 sg13g2_a21oi_1 _1621_ (.A1(_0708_),
    .A2(_0716_),
    .Y(_0010_),
    .B1(_0717_));
 sg13g2_nor4_1 _1622_ (.A(_0208_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0718_));
 sg13g2_nand4_1 _1623_ (.B(net299),
    .C(net297),
    .A(net351),
    .Y(_0719_),
    .D(_0588_));
 sg13g2_nand4_1 _1624_ (.B(net299),
    .C(net297),
    .A(net363),
    .Y(_0720_),
    .D(_0590_));
 sg13g2_a22oi_1 _1625_ (.Y(_0721_),
    .B1(_0593_),
    .B2(net342),
    .A2(_0592_),
    .A1(\u8.rc[26] ));
 sg13g2_nand4_1 _1626_ (.B(_0719_),
    .C(_0720_),
    .A(_0599_),
    .Y(_0722_),
    .D(_0721_));
 sg13g2_nand2_1 _1627_ (.Y(_0723_),
    .A(\u8.rc[26] ),
    .B(_0422_));
 sg13g2_nand3_1 _1628_ (.B(net312),
    .C(net311),
    .A(net342),
    .Y(_0724_));
 sg13g2_nand2_1 _1629_ (.Y(_0725_),
    .A(_0406_),
    .B(_0598_));
 sg13g2_a22oi_1 _1630_ (.Y(_0726_),
    .B1(_0427_),
    .B2(net363),
    .A2(_0426_),
    .A1(net351));
 sg13g2_a21oi_1 _1631_ (.A1(net373),
    .A2(_0604_),
    .Y(_0727_),
    .B1(_0725_));
 sg13g2_nand4_1 _1632_ (.B(_0724_),
    .C(_0726_),
    .A(_0723_),
    .Y(_0728_),
    .D(_0727_));
 sg13g2_nor2b_1 _1633_ (.A(_0603_),
    .B_N(_0728_),
    .Y(_0729_));
 sg13g2_o21ai_1 _1634_ (.B1(_0729_),
    .Y(_0730_),
    .A1(_0718_),
    .A2(_0722_));
 sg13g2_nor2_2 _1635_ (.A(\u8.ls[2] ),
    .B(net410),
    .Y(_0731_));
 sg13g2_inv_1 _1636_ (.Y(_0732_),
    .A(_0731_));
 sg13g2_nor3_1 _1637_ (.A(_0561_),
    .B(net329),
    .C(_0638_),
    .Y(_0733_));
 sg13g2_nor3_1 _1638_ (.A(net330),
    .B(_0625_),
    .C(_0731_),
    .Y(_0734_));
 sg13g2_o21ai_1 _1639_ (.B1(net306),
    .Y(_0735_),
    .A1(_0733_),
    .A2(_0734_));
 sg13g2_nor3_1 _1640_ (.A(_0497_),
    .B(_0619_),
    .C(_0638_),
    .Y(_0736_));
 sg13g2_a21oi_1 _1641_ (.A1(_0192_),
    .A2(net392),
    .Y(_0737_),
    .B1(_0625_));
 sg13g2_a221oi_1 _1642_ (.B2(net331),
    .C1(_0736_),
    .B1(_0737_),
    .A1(net373),
    .Y(_0738_),
    .A2(net327));
 sg13g2_nand2_2 _1643_ (.Y(_0739_),
    .A(\u8.hs[2] ),
    .B(net411));
 sg13g2_or2_1 _1644_ (.X(_0740_),
    .B(_0739_),
    .A(net329));
 sg13g2_a221oi_1 _1645_ (.B2(net327),
    .C1(net322),
    .B1(_0732_),
    .A1(_0562_),
    .Y(_0741_),
    .A2(_0632_));
 sg13g2_nand2_1 _1646_ (.Y(_0742_),
    .A(net356),
    .B(net392));
 sg13g2_a22oi_1 _1647_ (.Y(_0743_),
    .B1(_0742_),
    .B2(net322),
    .A2(_0741_),
    .A1(_0740_));
 sg13g2_a21oi_1 _1648_ (.A1(net320),
    .A2(_0743_),
    .Y(_0744_),
    .B1(_0476_));
 sg13g2_o21ai_1 _1649_ (.B1(_0744_),
    .Y(_0745_),
    .A1(net302),
    .A2(_0738_));
 sg13g2_nor2b_1 _1650_ (.A(_0745_),
    .B_N(_0735_),
    .Y(_0746_));
 sg13g2_o21ai_1 _1651_ (.B1(_0647_),
    .Y(_0747_),
    .A1(net373),
    .A2(net309));
 sg13g2_or3_1 _1652_ (.A(net301),
    .B(_0746_),
    .C(_0747_),
    .X(_0748_));
 sg13g2_a21o_1 _1653_ (.A2(_0748_),
    .A1(_0730_),
    .B1(net385),
    .X(_0749_));
 sg13g2_nor4_1 _1654_ (.A(\u8.rcop[1] ),
    .B(_0497_),
    .C(_0638_),
    .D(_0656_),
    .Y(_0750_));
 sg13g2_nor2_1 _1655_ (.A(\u8.rc[26] ),
    .B(net391),
    .Y(_0751_));
 sg13g2_nand2_1 _1656_ (.Y(_0752_),
    .A(net326),
    .B(_0732_));
 sg13g2_a21oi_1 _1657_ (.A1(_0215_),
    .A2(net391),
    .Y(_0753_),
    .B1(_0561_));
 sg13g2_a221oi_1 _1658_ (.B2(_0657_),
    .C1(_0750_),
    .B1(_0753_),
    .A1(_0663_),
    .Y(_0754_),
    .A2(_0737_));
 sg13g2_o21ai_1 _1659_ (.B1(_0754_),
    .Y(_0755_),
    .A1(_0751_),
    .A2(_0752_));
 sg13g2_a21oi_1 _1660_ (.A1(net336),
    .A2(_0755_),
    .Y(_0756_),
    .B1(_0652_));
 sg13g2_o21ai_1 _1661_ (.B1(net383),
    .Y(_0757_),
    .A1(net95),
    .A2(_0653_));
 sg13g2_a21oi_1 _1662_ (.A1(_0749_),
    .A2(_0756_),
    .Y(_0011_),
    .B1(_0757_));
 sg13g2_nor4_1 _1663_ (.A(_0207_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0758_));
 sg13g2_nand4_1 _1664_ (.B(net300),
    .C(net297),
    .A(net349),
    .Y(_0759_),
    .D(_0588_));
 sg13g2_nand4_1 _1665_ (.B(net300),
    .C(net297),
    .A(net362),
    .Y(_0760_),
    .D(_0590_));
 sg13g2_a22oi_1 _1666_ (.Y(_0761_),
    .B1(_0593_),
    .B2(net340),
    .A2(_0592_),
    .A1(net380));
 sg13g2_nand4_1 _1667_ (.B(_0759_),
    .C(_0760_),
    .A(_0599_),
    .Y(_0762_),
    .D(_0761_));
 sg13g2_nand2_1 _1668_ (.Y(_0763_),
    .A(\u8.ls[3] ),
    .B(_0604_));
 sg13g2_a21oi_1 _1669_ (.A1(net349),
    .A2(_0426_),
    .Y(_0764_),
    .B1(_0422_));
 sg13g2_a221oi_1 _1670_ (.B2(net340),
    .C1(_0725_),
    .B1(_0428_),
    .A1(net362),
    .Y(_0765_),
    .A2(_0427_));
 sg13g2_nand3_1 _1671_ (.B(_0764_),
    .C(_0765_),
    .A(_0763_),
    .Y(_0766_));
 sg13g2_nor2b_1 _1672_ (.A(_0603_),
    .B_N(_0766_),
    .Y(_0767_));
 sg13g2_o21ai_1 _1673_ (.B1(_0767_),
    .Y(_0768_),
    .A1(_0758_),
    .A2(_0762_));
 sg13g2_nor2_1 _1674_ (.A(\u8.ls[3] ),
    .B(net409),
    .Y(_0769_));
 sg13g2_nand2_1 _1675_ (.Y(_0770_),
    .A(_0207_),
    .B(net391));
 sg13g2_nor3_1 _1676_ (.A(net333),
    .B(_0691_),
    .C(_0769_),
    .Y(_0771_));
 sg13g2_nand2_1 _1677_ (.Y(_0772_),
    .A(_0567_),
    .B(net330));
 sg13g2_nor2_1 _1678_ (.A(_0699_),
    .B(_0772_),
    .Y(_0773_));
 sg13g2_o21ai_1 _1679_ (.B1(net306),
    .Y(_0774_),
    .A1(_0771_),
    .A2(_0773_));
 sg13g2_a21oi_1 _1680_ (.A1(_0191_),
    .A2(net406),
    .Y(_0775_),
    .B1(_0699_));
 sg13g2_o21ai_1 _1681_ (.B1(_0511_),
    .Y(_0776_),
    .A1(net357),
    .A2(net403));
 sg13g2_a21oi_1 _1682_ (.A1(_0191_),
    .A2(_0222_),
    .Y(_0777_),
    .B1(_0691_));
 sg13g2_a22oi_1 _1683_ (.Y(_0778_),
    .B1(_0777_),
    .B2(net331),
    .A2(net327),
    .A1(\u8.ls[3] ));
 sg13g2_o21ai_1 _1684_ (.B1(_0778_),
    .Y(_0779_),
    .A1(_0619_),
    .A2(_0776_));
 sg13g2_nand2_2 _1685_ (.Y(_0780_),
    .A(_0200_),
    .B(net394));
 sg13g2_nand2_1 _1686_ (.Y(_0781_),
    .A(net322),
    .B(_0780_));
 sg13g2_o21ai_1 _1687_ (.B1(net330),
    .Y(_0782_),
    .A1(net354),
    .A2(net391));
 sg13g2_a22oi_1 _1688_ (.Y(_0783_),
    .B1(_0770_),
    .B2(net327),
    .A2(_0632_),
    .A1(_0567_));
 sg13g2_nand3_1 _1689_ (.B(_0782_),
    .C(_0783_),
    .A(_0781_),
    .Y(_0784_));
 sg13g2_a221oi_1 _1690_ (.B2(net320),
    .C1(_0476_),
    .B1(_0784_),
    .A1(_0574_),
    .Y(_0785_),
    .A2(_0779_));
 sg13g2_a22oi_1 _1691_ (.Y(_0786_),
    .B1(_0774_),
    .B2(_0785_),
    .A2(_0476_),
    .A1(_0207_));
 sg13g2_nand2_1 _1692_ (.Y(_0787_),
    .A(_0684_),
    .B(_0786_));
 sg13g2_a21o_1 _1693_ (.A2(_0787_),
    .A1(_0768_),
    .B1(net385),
    .X(_0788_));
 sg13g2_nor2_1 _1694_ (.A(net380),
    .B(net391),
    .Y(_0789_));
 sg13g2_nand2_1 _1695_ (.Y(_0790_),
    .A(net326),
    .B(_0770_));
 sg13g2_o21ai_1 _1696_ (.B1(_0567_),
    .Y(_0791_),
    .A1(\u8.rc[27] ),
    .A2(net402));
 sg13g2_nor2_1 _1697_ (.A(_0658_),
    .B(_0791_),
    .Y(_0792_));
 sg13g2_a221oi_1 _1698_ (.B2(_0663_),
    .C1(_0792_),
    .B1(_0777_),
    .A1(_0661_),
    .Y(_0793_),
    .A2(_0775_));
 sg13g2_o21ai_1 _1699_ (.B1(_0793_),
    .Y(_0794_),
    .A1(_0789_),
    .A2(_0790_));
 sg13g2_a21oi_1 _1700_ (.A1(net336),
    .A2(_0794_),
    .Y(_0795_),
    .B1(_0652_));
 sg13g2_o21ai_1 _1701_ (.B1(net383),
    .Y(_0796_),
    .A1(net94),
    .A2(_0653_));
 sg13g2_a21oi_1 _1702_ (.A1(_0788_),
    .A2(_0795_),
    .Y(_0012_),
    .B1(_0796_));
 sg13g2_nor4_1 _1703_ (.A(_0206_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0797_));
 sg13g2_nand4_1 _1704_ (.B(net300),
    .C(net298),
    .A(net347),
    .Y(_0798_),
    .D(_0588_));
 sg13g2_nand4_1 _1705_ (.B(net300),
    .C(net298),
    .A(net359),
    .Y(_0799_),
    .D(_0590_));
 sg13g2_nand3_1 _1706_ (.B(\u8.rc[28] ),
    .C(_0592_),
    .A(_0212_),
    .Y(_0800_));
 sg13g2_a21oi_1 _1707_ (.A1(net339),
    .A2(_0593_),
    .Y(_0801_),
    .B1(_0598_));
 sg13g2_nand4_1 _1708_ (.B(_0799_),
    .C(_0800_),
    .A(_0798_),
    .Y(_0802_),
    .D(_0801_));
 sg13g2_and2_1 _1709_ (.A(net347),
    .B(_0426_),
    .X(_0803_));
 sg13g2_a21oi_1 _1710_ (.A1(net359),
    .A2(_0427_),
    .Y(_0804_),
    .B1(_0803_));
 sg13g2_nand3_1 _1711_ (.B(_0598_),
    .C(_0804_),
    .A(_0396_),
    .Y(_0805_));
 sg13g2_a21oi_1 _1712_ (.A1(net371),
    .A2(_0604_),
    .Y(_0806_),
    .B1(_0805_));
 sg13g2_nor2_1 _1713_ (.A(_0603_),
    .B(_0806_),
    .Y(_0807_));
 sg13g2_o21ai_1 _1714_ (.B1(_0807_),
    .Y(_0808_),
    .A1(_0797_),
    .A2(_0802_));
 sg13g2_nand2b_1 _1715_ (.Y(_0809_),
    .B(_0742_),
    .A_N(_0523_));
 sg13g2_nor2b_1 _1716_ (.A(_0619_),
    .B_N(_0809_),
    .Y(_0810_));
 sg13g2_o21ai_1 _1717_ (.B1(_0739_),
    .Y(_0811_),
    .A1(_0190_),
    .A2(net404));
 sg13g2_a221oi_1 _1718_ (.B2(net333),
    .C1(_0810_),
    .B1(_0811_),
    .A1(net371),
    .Y(_0812_),
    .A2(_0618_));
 sg13g2_nor2_1 _1719_ (.A(net351),
    .B(net403),
    .Y(_0813_));
 sg13g2_or2_1 _1720_ (.X(_0814_),
    .B(net405),
    .A(net351));
 sg13g2_nor2_2 _1721_ (.A(net372),
    .B(net410),
    .Y(_0815_));
 sg13g2_nor2b_1 _1722_ (.A(_0815_),
    .B_N(_0618_),
    .Y(_0816_));
 sg13g2_nand2b_2 _1723_ (.Y(_0817_),
    .B(net408),
    .A_N(net352));
 sg13g2_a221oi_1 _1724_ (.B2(net333),
    .C1(_0816_),
    .B1(_0817_),
    .A1(_0558_),
    .Y(_0818_),
    .A2(_0632_));
 sg13g2_o21ai_1 _1725_ (.B1(_0818_),
    .Y(_0819_),
    .A1(_0636_),
    .A2(_0813_));
 sg13g2_a21oi_1 _1726_ (.A1(net320),
    .A2(_0819_),
    .Y(_0820_),
    .B1(_0476_));
 sg13g2_o21ai_1 _1727_ (.B1(_0820_),
    .Y(_0821_),
    .A1(net302),
    .A2(_0812_));
 sg13g2_a21oi_1 _1728_ (.A1(_0201_),
    .A2(net404),
    .Y(_0822_),
    .B1(_0815_));
 sg13g2_and2_1 _1729_ (.A(_0557_),
    .B(_0742_),
    .X(_0823_));
 sg13g2_nor2_1 _1730_ (.A(net332),
    .B(_0822_),
    .Y(_0824_));
 sg13g2_a21oi_1 _1731_ (.A1(net332),
    .A2(_0823_),
    .Y(_0825_),
    .B1(_0824_));
 sg13g2_a21oi_1 _1732_ (.A1(net306),
    .A2(_0825_),
    .Y(_0826_),
    .B1(_0821_));
 sg13g2_o21ai_1 _1733_ (.B1(_0647_),
    .Y(_0827_),
    .A1(net371),
    .A2(net309));
 sg13g2_or3_1 _1734_ (.A(_0390_),
    .B(_0826_),
    .C(_0827_),
    .X(_0828_));
 sg13g2_a21o_1 _1735_ (.A2(_0828_),
    .A1(_0808_),
    .B1(net385),
    .X(_0829_));
 sg13g2_o21ai_1 _1736_ (.B1(_0557_),
    .Y(_0830_),
    .A1(_0214_),
    .A2(net404));
 sg13g2_a22oi_1 _1737_ (.Y(_0831_),
    .B1(_0830_),
    .B2(_0657_),
    .A2(_0811_),
    .A1(_0663_));
 sg13g2_a21oi_1 _1738_ (.A1(_0214_),
    .A2(net403),
    .Y(_0832_),
    .B1(_0815_));
 sg13g2_a22oi_1 _1739_ (.Y(_0833_),
    .B1(_0832_),
    .B2(_0660_),
    .A2(_0809_),
    .A1(_0661_));
 sg13g2_nand2_1 _1740_ (.Y(_0834_),
    .A(_0831_),
    .B(_0833_));
 sg13g2_a21oi_1 _1741_ (.A1(net336),
    .A2(_0834_),
    .Y(_0835_),
    .B1(_0652_));
 sg13g2_o21ai_1 _1742_ (.B1(net384),
    .Y(_0836_),
    .A1(net89),
    .A2(_0653_));
 sg13g2_a21oi_1 _1743_ (.A1(_0829_),
    .A2(_0835_),
    .Y(_0013_),
    .B1(_0836_));
 sg13g2_nor4_1 _1744_ (.A(_0205_),
    .B(_0589_),
    .C(_0591_),
    .D(_0594_),
    .Y(_0837_));
 sg13g2_nand4_1 _1745_ (.B(net299),
    .C(net298),
    .A(net346),
    .Y(_0838_),
    .D(_0588_));
 sg13g2_nand4_1 _1746_ (.B(net299),
    .C(net298),
    .A(net357),
    .Y(_0839_),
    .D(_0590_));
 sg13g2_nand3_1 _1747_ (.B(\u8.rc[29] ),
    .C(_0592_),
    .A(_0212_),
    .Y(_0840_));
 sg13g2_a21oi_1 _1748_ (.A1(net338),
    .A2(_0593_),
    .Y(_0841_),
    .B1(_0598_));
 sg13g2_nand4_1 _1749_ (.B(_0839_),
    .C(_0840_),
    .A(_0838_),
    .Y(_0842_),
    .D(_0841_));
 sg13g2_nand2_1 _1750_ (.Y(_0843_),
    .A(_0202_),
    .B(_0427_));
 sg13g2_o21ai_1 _1751_ (.B1(_0843_),
    .Y(_0844_),
    .A1(net370),
    .A2(_0605_));
 sg13g2_a21oi_1 _1752_ (.A1(_0598_),
    .A2(_0844_),
    .Y(_0845_),
    .B1(_0603_));
 sg13g2_o21ai_1 _1753_ (.B1(_0845_),
    .Y(_0846_),
    .A1(_0837_),
    .A2(_0842_));
 sg13g2_nand2_2 _1754_ (.Y(_0847_),
    .A(net350),
    .B(net407));
 sg13g2_nor2_1 _1755_ (.A(_0205_),
    .B(net392),
    .Y(_0848_));
 sg13g2_nor2_2 _1756_ (.A(_0205_),
    .B(net407),
    .Y(_0849_));
 sg13g2_nand2_1 _1757_ (.Y(_0850_),
    .A(net328),
    .B(_0849_));
 sg13g2_nor2_1 _1758_ (.A(_0199_),
    .B(net401),
    .Y(_0851_));
 sg13g2_o21ai_1 _1759_ (.B1(_0850_),
    .Y(_0852_),
    .A1(net329),
    .A2(_0847_));
 sg13g2_a221oi_1 _1760_ (.B2(net322),
    .C1(_0852_),
    .B1(_0851_),
    .A1(_0632_),
    .Y(_0853_),
    .A2(_0848_));
 sg13g2_o21ai_1 _1761_ (.B1(net309),
    .Y(_0854_),
    .A1(_0380_),
    .A2(_0853_));
 sg13g2_o21ai_1 _1762_ (.B1(_0780_),
    .Y(_0855_),
    .A1(net340),
    .A2(net391));
 sg13g2_nand2_2 _1763_ (.Y(_0856_),
    .A(net354),
    .B(net413));
 sg13g2_o21ai_1 _1764_ (.B1(_0856_),
    .Y(_0857_),
    .A1(_0189_),
    .A2(net405));
 sg13g2_a22oi_1 _1765_ (.Y(_0858_),
    .B1(_0857_),
    .B2(net330),
    .A2(net327),
    .A1(net370));
 sg13g2_o21ai_1 _1766_ (.B1(_0858_),
    .Y(_0859_),
    .A1(_0619_),
    .A2(_0855_));
 sg13g2_nor2b_1 _1767_ (.A(_0849_),
    .B_N(_0856_),
    .Y(_0860_));
 sg13g2_a21o_1 _1768_ (.A2(_0780_),
    .A1(_0555_),
    .B1(net329),
    .X(_0861_));
 sg13g2_a21oi_1 _1769_ (.A1(net329),
    .A2(_0860_),
    .Y(_0862_),
    .B1(net303));
 sg13g2_a221oi_1 _1770_ (.B2(_0862_),
    .C1(_0854_),
    .B1(_0861_),
    .A1(_0574_),
    .Y(_0863_),
    .A2(_0859_));
 sg13g2_o21ai_1 _1771_ (.B1(_0647_),
    .Y(_0864_),
    .A1(net370),
    .A2(net309));
 sg13g2_or3_1 _1772_ (.A(net301),
    .B(_0863_),
    .C(_0864_),
    .X(_0865_));
 sg13g2_a21o_1 _1773_ (.A2(_0865_),
    .A1(_0846_),
    .B1(_0584_),
    .X(_0866_));
 sg13g2_nor3_1 _1774_ (.A(\u8.rcop[1] ),
    .B(_0656_),
    .C(_0855_),
    .Y(_0867_));
 sg13g2_nor2_1 _1775_ (.A(net326),
    .B(_0867_),
    .Y(_0868_));
 sg13g2_mux2_1 _1776_ (.A0(\u8.rc[29] ),
    .A1(net370),
    .S(net400),
    .X(_0869_));
 sg13g2_a22oi_1 _1777_ (.Y(_0870_),
    .B1(_0869_),
    .B2(_0657_),
    .A2(_0857_),
    .A1(_0663_));
 sg13g2_a21oi_1 _1778_ (.A1(net132),
    .A2(net400),
    .Y(_0871_),
    .B1(_0849_));
 sg13g2_a22oi_1 _1779_ (.Y(_0872_),
    .B1(_0871_),
    .B2(net326),
    .A2(_0870_),
    .A1(_0868_));
 sg13g2_a21oi_1 _1780_ (.A1(_0665_),
    .A2(_0872_),
    .Y(_0873_),
    .B1(_0652_));
 sg13g2_o21ai_1 _1781_ (.B1(net384),
    .Y(_0874_),
    .A1(net93),
    .A2(_0653_));
 sg13g2_a21oi_1 _1782_ (.A1(_0866_),
    .A2(_0873_),
    .Y(_0014_),
    .B1(_0874_));
 sg13g2_o21ai_1 _1783_ (.B1(_0598_),
    .Y(_0875_),
    .A1(net368),
    .A2(_0605_));
 sg13g2_nor2_1 _1784_ (.A(\u8.ls[6] ),
    .B(net408),
    .Y(_0876_));
 sg13g2_o21ai_1 _1785_ (.B1(_0817_),
    .Y(_0877_),
    .A1(net369),
    .A2(net405));
 sg13g2_a21oi_1 _1786_ (.A1(_0565_),
    .A2(_0814_),
    .Y(_0878_),
    .B1(net329));
 sg13g2_a21oi_1 _1787_ (.A1(_0616_),
    .A2(_0877_),
    .Y(_0879_),
    .B1(_0878_));
 sg13g2_nor3_1 _1788_ (.A(_0538_),
    .B(_0619_),
    .C(_0813_),
    .Y(_0880_));
 sg13g2_mux2_1 _1789_ (.A0(net339),
    .A1(net351),
    .S(net401),
    .X(_0881_));
 sg13g2_a221oi_1 _1790_ (.B2(net333),
    .C1(_0880_),
    .B1(_0881_),
    .A1(net368),
    .Y(_0882_),
    .A2(net328));
 sg13g2_nand2_1 _1791_ (.Y(_0883_),
    .A(net348),
    .B(net405));
 sg13g2_nand2b_1 _1792_ (.Y(_0884_),
    .B(net328),
    .A_N(_0876_));
 sg13g2_a221oi_1 _1793_ (.B2(net333),
    .C1(_0635_),
    .B1(_0883_),
    .A1(_0565_),
    .Y(_0885_),
    .A2(_0632_));
 sg13g2_a22oi_1 _1794_ (.Y(_0886_),
    .B1(_0884_),
    .B2(_0885_),
    .A2(net322),
    .A1(_0621_));
 sg13g2_nand2_1 _1795_ (.Y(_0887_),
    .A(net320),
    .B(_0886_));
 sg13g2_o21ai_1 _1796_ (.B1(_0887_),
    .Y(_0888_),
    .A1(net302),
    .A2(_0882_));
 sg13g2_a221oi_1 _1797_ (.B2(net306),
    .C1(_0888_),
    .B1(_0879_),
    .A1(net368),
    .Y(_0889_),
    .A2(_0476_));
 sg13g2_nand2b_1 _1798_ (.Y(_0890_),
    .B(_0684_),
    .A_N(_0889_));
 sg13g2_o21ai_1 _1799_ (.B1(_0890_),
    .Y(_0891_),
    .A1(_0603_),
    .A2(_0875_));
 sg13g2_nand2_1 _1800_ (.Y(_0892_),
    .A(_0213_),
    .B(net392));
 sg13g2_nand3_1 _1801_ (.B(_0657_),
    .C(_0892_),
    .A(_0565_),
    .Y(_0893_));
 sg13g2_nand3b_1 _1802_ (.B(_0661_),
    .C(_0814_),
    .Y(_0894_),
    .A_N(_0538_));
 sg13g2_a21oi_1 _1803_ (.A1(_0213_),
    .A2(net405),
    .Y(_0895_),
    .B1(_0876_));
 sg13g2_a22oi_1 _1804_ (.Y(_0896_),
    .B1(_0895_),
    .B2(net326),
    .A2(_0881_),
    .A1(_0663_));
 sg13g2_nand3_1 _1805_ (.B(_0894_),
    .C(_0896_),
    .A(_0893_),
    .Y(_0897_));
 sg13g2_a221oi_1 _1806_ (.B2(net336),
    .C1(_0652_),
    .B1(_0897_),
    .A1(_0585_),
    .Y(_0898_),
    .A2(_0891_));
 sg13g2_o21ai_1 _1807_ (.B1(net383),
    .Y(_0899_),
    .A1(net86),
    .A2(_0653_));
 sg13g2_nor2_1 _1808_ (.A(_0898_),
    .B(_0899_),
    .Y(_0015_));
 sg13g2_a21oi_1 _1809_ (.A1(_0287_),
    .A2(_0288_),
    .Y(_0900_),
    .B1(_0603_));
 sg13g2_nor3_1 _1810_ (.A(_0552_),
    .B(net329),
    .C(_0851_),
    .Y(_0901_));
 sg13g2_nor2_1 _1811_ (.A(net367),
    .B(net408),
    .Y(_0902_));
 sg13g2_or2_1 _1812_ (.X(_0903_),
    .B(net400),
    .A(net365));
 sg13g2_nand2_1 _1813_ (.Y(_0904_),
    .A(_0199_),
    .B(net401));
 sg13g2_a21oi_1 _1814_ (.A1(_0903_),
    .A2(_0904_),
    .Y(_0905_),
    .B1(net330));
 sg13g2_nor3_1 _1815_ (.A(net303),
    .B(_0901_),
    .C(_0905_),
    .Y(_0906_));
 sg13g2_nand2b_1 _1816_ (.Y(_0907_),
    .B(_0276_),
    .A_N(_0238_));
 sg13g2_o21ai_1 _1817_ (.B1(net322),
    .Y(_0908_),
    .A1(net400),
    .A2(_0907_));
 sg13g2_a22oi_1 _1818_ (.Y(_0909_),
    .B1(_0903_),
    .B2(net327),
    .A2(_0632_),
    .A1(_0553_));
 sg13g2_o21ai_1 _1819_ (.B1(net330),
    .Y(_0910_),
    .A1(net391),
    .A2(_0907_));
 sg13g2_nand3_1 _1820_ (.B(_0909_),
    .C(_0910_),
    .A(_0908_),
    .Y(_0911_));
 sg13g2_and2_1 _1821_ (.A(net320),
    .B(_0911_),
    .X(_0912_));
 sg13g2_a21oi_1 _1822_ (.A1(net338),
    .A2(net401),
    .Y(_0913_),
    .B1(_0851_));
 sg13g2_o21ai_1 _1823_ (.B1(_0847_),
    .Y(_0914_),
    .A1(_0188_),
    .A2(net407));
 sg13g2_a22oi_1 _1824_ (.Y(_0915_),
    .B1(_0914_),
    .B2(net330),
    .A2(net327),
    .A1(net365));
 sg13g2_o21ai_1 _1825_ (.B1(_0915_),
    .Y(_0916_),
    .A1(_0619_),
    .A2(_0913_));
 sg13g2_nor2b_1 _1826_ (.A(net302),
    .B_N(_0916_),
    .Y(_0917_));
 sg13g2_nor4_1 _1827_ (.A(_0476_),
    .B(_0906_),
    .C(_0912_),
    .D(_0917_),
    .Y(_0918_));
 sg13g2_o21ai_1 _1828_ (.B1(_0647_),
    .Y(_0919_),
    .A1(net365),
    .A2(net309));
 sg13g2_nor3_1 _1829_ (.A(net301),
    .B(_0918_),
    .C(_0919_),
    .Y(_0920_));
 sg13g2_o21ai_1 _1830_ (.B1(_0585_),
    .Y(_0921_),
    .A1(_0900_),
    .A2(_0920_));
 sg13g2_nor2_1 _1831_ (.A(_0212_),
    .B(net401),
    .Y(_0922_));
 sg13g2_o21ai_1 _1832_ (.B1(_0657_),
    .Y(_0923_),
    .A1(_0552_),
    .A2(_0922_));
 sg13g2_nand2b_1 _1833_ (.Y(_0924_),
    .B(_0661_),
    .A_N(_0913_));
 sg13g2_a21oi_1 _1834_ (.A1(_0212_),
    .A2(net401),
    .Y(_0925_),
    .B1(_0902_));
 sg13g2_a22oi_1 _1835_ (.Y(_0926_),
    .B1(_0925_),
    .B2(net326),
    .A2(_0914_),
    .A1(_0663_));
 sg13g2_nand3_1 _1836_ (.B(_0924_),
    .C(_0926_),
    .A(_0923_),
    .Y(_0927_));
 sg13g2_a21oi_1 _1837_ (.A1(_0665_),
    .A2(_0927_),
    .Y(_0928_),
    .B1(_0652_));
 sg13g2_o21ai_1 _1838_ (.B1(net384),
    .Y(_0929_),
    .A1(net91),
    .A2(_0653_));
 sg13g2_a21oi_1 _1839_ (.A1(_0921_),
    .A2(_0928_),
    .Y(_0016_),
    .B1(_0929_));
 sg13g2_nor2_1 _1840_ (.A(\u8.rcip[2] ),
    .B(\u8.rcip[0] ),
    .Y(_0930_));
 sg13g2_nor3_2 _1841_ (.A(\u8.rcip[2] ),
    .B(\u8.rcip[1] ),
    .C(\u8.rcip[0] ),
    .Y(_0931_));
 sg13g2_nand2_1 _1842_ (.Y(_0932_),
    .A(_0197_),
    .B(_0930_));
 sg13g2_nor2_2 _1843_ (.A(_0459_),
    .B(_0478_),
    .Y(_0933_));
 sg13g2_a221oi_1 _1844_ (.B2(_0460_),
    .C1(_0461_),
    .B1(_0933_),
    .A1(net390),
    .Y(_0934_),
    .A2(_0932_));
 sg13g2_o21ai_1 _1845_ (.B1(net421),
    .Y(_0017_),
    .A1(_0211_),
    .A2(_0934_));
 sg13g2_nand2_1 _1846_ (.Y(_0935_),
    .A(net393),
    .B(net323));
 sg13g2_nor2b_2 _1847_ (.A(_0470_),
    .B_N(_0935_),
    .Y(_0936_));
 sg13g2_nand2b_2 _1848_ (.Y(_0937_),
    .B(_0935_),
    .A_N(_0470_));
 sg13g2_nor3_2 _1849_ (.A(\u8.rcip[2] ),
    .B(_0197_),
    .C(net413),
    .Y(_0938_));
 sg13g2_and2_1 _1850_ (.A(_0198_),
    .B(_0938_),
    .X(_0939_));
 sg13g2_a21oi_2 _1851_ (.B1(_0937_),
    .Y(_0940_),
    .A2(_0939_),
    .A1(net387));
 sg13g2_a21o_1 _1852_ (.A2(net8),
    .A1(net409),
    .B1(_0628_),
    .X(_0941_));
 sg13g2_nor2_2 _1853_ (.A(_0931_),
    .B(_0938_),
    .Y(_0942_));
 sg13g2_a22oi_1 _1854_ (.Y(_0943_),
    .B1(_0941_),
    .B2(_0942_),
    .A2(_0931_),
    .A1(net8));
 sg13g2_nor2_1 _1855_ (.A(_0445_),
    .B(_0478_),
    .Y(_0944_));
 sg13g2_nand2_2 _1856_ (.Y(_0945_),
    .A(net303),
    .B(net295));
 sg13g2_nand2_1 _1857_ (.Y(_0946_),
    .A(_0383_),
    .B(_0576_));
 sg13g2_nor2_2 _1858_ (.A(_0571_),
    .B(_0573_),
    .Y(_0947_));
 sg13g2_a22oi_1 _1859_ (.Y(_0948_),
    .B1(net292),
    .B2(net364),
    .A2(net293),
    .A1(_0941_));
 sg13g2_inv_1 _1860_ (.Y(_0949_),
    .A(_0948_));
 sg13g2_a221oi_1 _1861_ (.B2(net295),
    .C1(net388),
    .B1(_0949_),
    .A1(net8),
    .Y(_0950_),
    .A2(_0945_));
 sg13g2_a21o_1 _1862_ (.A2(_0943_),
    .A1(net388),
    .B1(_0950_),
    .X(_0951_));
 sg13g2_o21ai_1 _1863_ (.B1(net420),
    .Y(_0952_),
    .A1(net108),
    .A2(net289));
 sg13g2_a21oi_1 _1864_ (.A1(net289),
    .A2(_0951_),
    .Y(_0018_),
    .B1(_0952_));
 sg13g2_a21oi_1 _1865_ (.A1(net412),
    .A2(_0227_),
    .Y(_0953_),
    .B1(_0693_));
 sg13g2_a22oi_1 _1866_ (.Y(_0954_),
    .B1(_0942_),
    .B2(_0953_),
    .A2(_0931_),
    .A1(net9));
 sg13g2_a22oi_1 _1867_ (.Y(_0955_),
    .B1(_0953_),
    .B2(net293),
    .A2(net292),
    .A1(net361));
 sg13g2_inv_1 _1868_ (.Y(_0956_),
    .A(_0955_));
 sg13g2_a221oi_1 _1869_ (.B2(net295),
    .C1(net388),
    .B1(_0956_),
    .A1(net9),
    .Y(_0957_),
    .A2(_0945_));
 sg13g2_a21o_1 _1870_ (.A2(_0954_),
    .A1(net388),
    .B1(_0957_),
    .X(_0958_));
 sg13g2_o21ai_1 _1871_ (.B1(net420),
    .Y(_0959_),
    .A1(net374),
    .A2(net289));
 sg13g2_a21oi_1 _1872_ (.A1(net289),
    .A2(_0958_),
    .Y(_0019_),
    .B1(_0959_));
 sg13g2_a21oi_1 _1873_ (.A1(_0221_),
    .A2(net412),
    .Y(_0960_),
    .B1(_0731_));
 sg13g2_a22oi_1 _1874_ (.Y(_0961_),
    .B1(_0942_),
    .B2(_0960_),
    .A2(_0931_),
    .A1(net10));
 sg13g2_a22oi_1 _1875_ (.Y(_0962_),
    .B1(_0960_),
    .B2(net293),
    .A2(net292),
    .A1(net360));
 sg13g2_inv_1 _1876_ (.Y(_0963_),
    .A(_0962_));
 sg13g2_a221oi_1 _1877_ (.B2(net295),
    .C1(net388),
    .B1(_0963_),
    .A1(net10),
    .Y(_0964_),
    .A2(_0945_));
 sg13g2_a21o_1 _1878_ (.A2(_0961_),
    .A1(net390),
    .B1(_0964_),
    .X(_0965_));
 sg13g2_o21ai_1 _1879_ (.B1(net419),
    .Y(_0966_),
    .A1(net101),
    .A2(net288));
 sg13g2_a21oi_1 _1880_ (.A1(net288),
    .A2(_0965_),
    .Y(_0020_),
    .B1(_0966_));
 sg13g2_a21oi_1 _1881_ (.A1(net412),
    .A2(_0223_),
    .Y(_0967_),
    .B1(_0769_));
 sg13g2_a22oi_1 _1882_ (.Y(_0968_),
    .B1(_0942_),
    .B2(_0967_),
    .A2(_0931_),
    .A1(net11));
 sg13g2_a22oi_1 _1883_ (.Y(_0969_),
    .B1(_0967_),
    .B2(net293),
    .A2(_0947_),
    .A1(net358));
 sg13g2_inv_1 _1884_ (.Y(_0970_),
    .A(_0969_));
 sg13g2_a221oi_1 _1885_ (.B2(net296),
    .C1(net389),
    .B1(_0970_),
    .A1(net11),
    .Y(_0971_),
    .A2(_0945_));
 sg13g2_a21o_1 _1886_ (.A2(_0968_),
    .A1(net389),
    .B1(_0971_),
    .X(_0972_));
 sg13g2_o21ai_1 _1887_ (.B1(net420),
    .Y(_0973_),
    .A1(net109),
    .A2(net288));
 sg13g2_a21oi_1 _1888_ (.A1(net288),
    .A2(_0972_),
    .Y(_0021_),
    .B1(_0973_));
 sg13g2_a21oi_1 _1889_ (.A1(net410),
    .A2(_0224_),
    .Y(_0974_),
    .B1(_0815_));
 sg13g2_a22oi_1 _1890_ (.Y(_0975_),
    .B1(_0942_),
    .B2(_0974_),
    .A2(_0931_),
    .A1(net12));
 sg13g2_a22oi_1 _1891_ (.Y(_0976_),
    .B1(_0974_),
    .B2(net293),
    .A2(_0947_),
    .A1(net356));
 sg13g2_inv_1 _1892_ (.Y(_0977_),
    .A(_0976_));
 sg13g2_a221oi_1 _1893_ (.B2(net295),
    .C1(net388),
    .B1(_0977_),
    .A1(net12),
    .Y(_0978_),
    .A2(_0945_));
 sg13g2_a21o_1 _1894_ (.A2(_0975_),
    .A1(net389),
    .B1(_0978_),
    .X(_0979_));
 sg13g2_o21ai_1 _1895_ (.B1(net420),
    .Y(_0980_),
    .A1(net371),
    .A2(net289));
 sg13g2_a21oi_1 _1896_ (.A1(_0940_),
    .A2(_0979_),
    .Y(_0022_),
    .B1(_0980_));
 sg13g2_a21o_1 _1897_ (.A2(net13),
    .A1(net412),
    .B1(_0849_),
    .X(_0981_));
 sg13g2_a22oi_1 _1898_ (.Y(_0982_),
    .B1(_0942_),
    .B2(_0981_),
    .A2(_0931_),
    .A1(net13));
 sg13g2_a22oi_1 _1899_ (.Y(_0983_),
    .B1(_0981_),
    .B2(_0946_),
    .A2(_0947_),
    .A1(net354));
 sg13g2_inv_1 _1900_ (.Y(_0984_),
    .A(_0983_));
 sg13g2_a221oi_1 _1901_ (.B2(net295),
    .C1(net388),
    .B1(_0984_),
    .A1(net13),
    .Y(_0985_),
    .A2(_0945_));
 sg13g2_a21o_1 _1902_ (.A2(_0982_),
    .A1(net388),
    .B1(_0985_),
    .X(_0986_));
 sg13g2_o21ai_1 _1903_ (.B1(net420),
    .Y(_0987_),
    .A1(net104),
    .A2(net289));
 sg13g2_a21oi_1 _1904_ (.A1(net289),
    .A2(_0986_),
    .Y(_0023_),
    .B1(_0987_));
 sg13g2_o21ai_1 _1905_ (.B1(_0479_),
    .Y(_0988_),
    .A1(_0450_),
    .A2(_0932_));
 sg13g2_o21ai_1 _1906_ (.B1(net14),
    .Y(_0989_),
    .A1(_0551_),
    .A2(_0988_));
 sg13g2_a21oi_1 _1907_ (.A1(_0219_),
    .A2(net409),
    .Y(_0990_),
    .B1(_0876_));
 sg13g2_a22oi_1 _1908_ (.Y(_0991_),
    .B1(_0990_),
    .B2(net293),
    .A2(net292),
    .A1(net352));
 sg13g2_nand2b_1 _1909_ (.Y(_0992_),
    .B(_0933_),
    .A_N(_0991_));
 sg13g2_nor3_2 _1910_ (.A(_0450_),
    .B(_0931_),
    .C(_0938_),
    .Y(_0993_));
 sg13g2_a22oi_1 _1911_ (.Y(_0994_),
    .B1(_0990_),
    .B2(net321),
    .A2(_0448_),
    .A1(\u8.ls[0] ));
 sg13g2_nand4_1 _1912_ (.B(_0989_),
    .C(_0992_),
    .A(net287),
    .Y(_0995_),
    .D(_0994_));
 sg13g2_o21ai_1 _1913_ (.B1(net419),
    .Y(_0996_),
    .A1(net369),
    .A2(net286));
 sg13g2_nor2b_1 _1914_ (.A(_0996_),
    .B_N(_0995_),
    .Y(_0024_));
 sg13g2_nand2_1 _1915_ (.Y(_0997_),
    .A(net15),
    .B(_0988_));
 sg13g2_a21oi_1 _1916_ (.A1(_0220_),
    .A2(net414),
    .Y(_0998_),
    .B1(_0902_));
 sg13g2_a22oi_1 _1917_ (.Y(_0999_),
    .B1(_0998_),
    .B2(net293),
    .A2(net292),
    .A1(net350));
 sg13g2_inv_1 _1918_ (.Y(_1000_),
    .A(_0999_));
 sg13g2_o21ai_1 _1919_ (.B1(net315),
    .Y(_1001_),
    .A1(net374),
    .A2(net324));
 sg13g2_a22oi_1 _1920_ (.Y(_1002_),
    .B1(_1000_),
    .B2(_0933_),
    .A2(_0998_),
    .A1(net321));
 sg13g2_nand4_1 _1921_ (.B(_0997_),
    .C(_1001_),
    .A(net287),
    .Y(_1003_),
    .D(_1002_));
 sg13g2_o21ai_1 _1922_ (.B1(net417),
    .Y(_1004_),
    .A1(net367),
    .A2(net285));
 sg13g2_nor2b_1 _1923_ (.A(_1004_),
    .B_N(_1003_),
    .Y(_0025_));
 sg13g2_a21oi_1 _1924_ (.A1(net393),
    .A2(_0226_),
    .Y(_1005_),
    .B1(_0631_));
 sg13g2_a21oi_1 _1925_ (.A1(_0383_),
    .A2(_0576_),
    .Y(_1006_),
    .B1(_1005_));
 sg13g2_a221oi_1 _1926_ (.B2(_0194_),
    .C1(_1006_),
    .B1(net292),
    .A1(_0210_),
    .Y(_1007_),
    .A2(net305));
 sg13g2_nand2b_1 _1927_ (.Y(_1008_),
    .B(net295),
    .A_N(_1007_));
 sg13g2_nand2_1 _1928_ (.Y(_1009_),
    .A(net15),
    .B(net324));
 sg13g2_and2_1 _1929_ (.A(_0445_),
    .B(_1009_),
    .X(_1010_));
 sg13g2_nand2_1 _1930_ (.Y(_1011_),
    .A(_0445_),
    .B(_1009_));
 sg13g2_nand2_1 _1931_ (.Y(_1012_),
    .A(net101),
    .B(net334));
 sg13g2_a21oi_1 _1932_ (.A1(net310),
    .A2(_1012_),
    .Y(_1013_),
    .B1(net386));
 sg13g2_a22oi_1 _1933_ (.Y(_1014_),
    .B1(_1008_),
    .B2(_1013_),
    .A2(_1005_),
    .A1(net321));
 sg13g2_o21ai_1 _1934_ (.B1(net419),
    .Y(_1015_),
    .A1(net364),
    .A2(net288));
 sg13g2_a21oi_1 _1935_ (.A1(net288),
    .A2(_1014_),
    .Y(_0026_),
    .B1(_1015_));
 sg13g2_nand2_1 _1936_ (.Y(_1016_),
    .A(_0489_),
    .B(_0695_));
 sg13g2_nand2_1 _1937_ (.Y(_1017_),
    .A(net293),
    .B(_1016_));
 sg13g2_a22oi_1 _1938_ (.Y(_1018_),
    .B1(net292),
    .B2(_0193_),
    .A2(net304),
    .A1(_0209_));
 sg13g2_nand3_1 _1939_ (.B(_1017_),
    .C(_1018_),
    .A(_0933_),
    .Y(_0054_));
 sg13g2_o21ai_1 _1940_ (.B1(net315),
    .Y(_0055_),
    .A1(\u8.ls[3] ),
    .A2(net324));
 sg13g2_nand3_1 _1941_ (.B(_0695_),
    .C(net321),
    .A(_0489_),
    .Y(_0056_));
 sg13g2_nand4_1 _1942_ (.B(_0054_),
    .C(_0055_),
    .A(net287),
    .Y(_0057_),
    .D(_0056_));
 sg13g2_o21ai_1 _1943_ (.B1(net418),
    .Y(_0058_),
    .A1(net361),
    .A2(net285));
 sg13g2_nor2b_1 _1944_ (.A(_0058_),
    .B_N(_0057_),
    .Y(_0027_));
 sg13g2_nor2_1 _1945_ (.A(net373),
    .B(net303),
    .Y(_0059_));
 sg13g2_a21oi_1 _1946_ (.A1(net313),
    .A2(_0563_),
    .Y(_0060_),
    .B1(net292));
 sg13g2_o21ai_1 _1947_ (.B1(_0060_),
    .Y(_0061_),
    .A1(\u8.ls[8] ),
    .A2(_0576_));
 sg13g2_o21ai_1 _1948_ (.B1(net295),
    .Y(_0062_),
    .A1(_0059_),
    .A2(_0061_));
 sg13g2_nand2_1 _1949_ (.Y(_0063_),
    .A(net372),
    .B(net334));
 sg13g2_a21oi_1 _1950_ (.A1(net310),
    .A2(_0063_),
    .Y(_0064_),
    .B1(net387));
 sg13g2_a22oi_1 _1951_ (.Y(_0065_),
    .B1(_0062_),
    .B2(_0064_),
    .A2(net321),
    .A1(_0564_));
 sg13g2_o21ai_1 _1952_ (.B1(net419),
    .Y(_0066_),
    .A1(net360),
    .A2(net286));
 sg13g2_a21oi_1 _1953_ (.A1(net286),
    .A2(_0065_),
    .Y(_0028_),
    .B1(_0066_));
 sg13g2_a22oi_1 _1954_ (.Y(_0067_),
    .B1(_0569_),
    .B2(net313),
    .A2(net304),
    .A1(_0207_));
 sg13g2_o21ai_1 _1955_ (.B1(_0067_),
    .Y(_0068_),
    .A1(net361),
    .A2(_0576_));
 sg13g2_o21ai_1 _1956_ (.B1(_1010_),
    .Y(_0069_),
    .A1(_0205_),
    .A2(net325));
 sg13g2_a21oi_1 _1957_ (.A1(net294),
    .A2(_0068_),
    .Y(_0070_),
    .B1(net387));
 sg13g2_a22oi_1 _1958_ (.Y(_0071_),
    .B1(_0069_),
    .B2(_0070_),
    .A2(net321),
    .A1(_0568_));
 sg13g2_o21ai_1 _1959_ (.B1(net419),
    .Y(_0072_),
    .A1(net358),
    .A2(net286));
 sg13g2_a21oi_1 _1960_ (.A1(net286),
    .A2(_0071_),
    .Y(_0029_),
    .B1(_0072_));
 sg13g2_a22oi_1 _1961_ (.Y(_0073_),
    .B1(_0575_),
    .B2(_0203_),
    .A2(_0559_),
    .A1(net313));
 sg13g2_o21ai_1 _1962_ (.B1(_0073_),
    .Y(_0074_),
    .A1(net372),
    .A2(net303));
 sg13g2_nand3_1 _1963_ (.B(net334),
    .C(net316),
    .A(net369),
    .Y(_0075_));
 sg13g2_a22oi_1 _1964_ (.Y(_0076_),
    .B1(_0075_),
    .B2(net310),
    .A2(_0074_),
    .A1(net294));
 sg13g2_a22oi_1 _1965_ (.Y(_0077_),
    .B1(_0076_),
    .B2(_0450_),
    .A2(net321),
    .A1(_0560_));
 sg13g2_o21ai_1 _1966_ (.B1(net420),
    .Y(_0078_),
    .A1(net103),
    .A2(net288));
 sg13g2_a21oi_1 _1967_ (.A1(net288),
    .A2(_0077_),
    .Y(_0030_),
    .B1(_0078_));
 sg13g2_nand2b_1 _1968_ (.Y(_0079_),
    .B(net321),
    .A_N(_0556_));
 sg13g2_a21oi_1 _1969_ (.A1(net367),
    .A2(net316),
    .Y(_0080_),
    .B1(net325));
 sg13g2_o21ai_1 _1970_ (.B1(_0079_),
    .Y(_0081_),
    .A1(_0451_),
    .A2(_0080_));
 sg13g2_a21oi_1 _1971_ (.A1(net357),
    .A2(_0571_),
    .Y(_0082_),
    .B1(_0573_));
 sg13g2_a221oi_1 _1972_ (.B2(net313),
    .C1(_0082_),
    .B1(_0556_),
    .A1(_0205_),
    .Y(_0083_),
    .A2(net304));
 sg13g2_a21oi_1 _1973_ (.A1(_0933_),
    .A2(_0083_),
    .Y(_0084_),
    .B1(_0081_));
 sg13g2_o21ai_1 _1974_ (.B1(net418),
    .Y(_0085_),
    .A1(net355),
    .A2(net285));
 sg13g2_a21oi_1 _1975_ (.A1(net285),
    .A2(_0084_),
    .Y(_0031_),
    .B1(_0085_));
 sg13g2_nor2_1 _1976_ (.A(net369),
    .B(net303),
    .Y(_0086_));
 sg13g2_nand2_1 _1977_ (.Y(_0087_),
    .A(_0201_),
    .B(_0575_));
 sg13g2_o21ai_1 _1978_ (.B1(_0087_),
    .Y(_0088_),
    .A1(_0383_),
    .A2(_0566_));
 sg13g2_o21ai_1 _1979_ (.B1(net294),
    .Y(_0089_),
    .A1(_0086_),
    .A2(_0088_));
 sg13g2_nand3_1 _1980_ (.B(net334),
    .C(net317),
    .A(net364),
    .Y(_0090_));
 sg13g2_a21oi_1 _1981_ (.A1(net310),
    .A2(_0090_),
    .Y(_0091_),
    .B1(net386));
 sg13g2_a22oi_1 _1982_ (.Y(_0092_),
    .B1(_0089_),
    .B2(_0091_),
    .A2(_0993_),
    .A1(_0566_));
 sg13g2_o21ai_1 _1983_ (.B1(net418),
    .Y(_0093_),
    .A1(net352),
    .A2(net285));
 sg13g2_a21oi_1 _1984_ (.A1(net285),
    .A2(_0092_),
    .Y(_0032_),
    .B1(_0093_));
 sg13g2_nor2_1 _1985_ (.A(net367),
    .B(net303),
    .Y(_0094_));
 sg13g2_nand2_1 _1986_ (.Y(_0095_),
    .A(_0200_),
    .B(_0575_));
 sg13g2_o21ai_1 _1987_ (.B1(_0095_),
    .Y(_0096_),
    .A1(_0383_),
    .A2(_0554_));
 sg13g2_o21ai_1 _1988_ (.B1(net296),
    .Y(_0097_),
    .A1(_0094_),
    .A2(_0096_));
 sg13g2_nand3_1 _1989_ (.B(net334),
    .C(net317),
    .A(net361),
    .Y(_0098_));
 sg13g2_a21oi_1 _1990_ (.A1(net310),
    .A2(_0098_),
    .Y(_0099_),
    .B1(net386));
 sg13g2_a22oi_1 _1991_ (.Y(_0100_),
    .B1(_0097_),
    .B2(_0099_),
    .A2(_0993_),
    .A1(_0554_));
 sg13g2_o21ai_1 _1992_ (.B1(net418),
    .Y(_0101_),
    .A1(net350),
    .A2(net285));
 sg13g2_a21oi_1 _1993_ (.A1(net285),
    .A2(_0100_),
    .Y(_0033_),
    .B1(_0101_));
 sg13g2_a21oi_1 _1994_ (.A1(net1),
    .A2(_0471_),
    .Y(_0102_),
    .B1(net75));
 sg13g2_nand3_1 _1995_ (.B(net1),
    .C(_0471_),
    .A(net75),
    .Y(_0103_));
 sg13g2_nand2_1 _1996_ (.Y(_0104_),
    .A(net419),
    .B(_0103_));
 sg13g2_nor2_1 _1997_ (.A(net76),
    .B(_0104_),
    .Y(_0034_));
 sg13g2_o21ai_1 _1998_ (.B1(net419),
    .Y(_0105_),
    .A1(_0197_),
    .A2(_0103_));
 sg13g2_a21oi_1 _1999_ (.A1(_0197_),
    .A2(_0103_),
    .Y(_0035_),
    .B1(_0105_));
 sg13g2_a21oi_1 _2000_ (.A1(net1),
    .A2(net323),
    .Y(_0106_),
    .B1(net84));
 sg13g2_nor2b_1 _2001_ (.A(_0106_),
    .B_N(net419),
    .Y(_0036_));
 sg13g2_o21ai_1 _2002_ (.B1(net383),
    .Y(_0107_),
    .A1(net70),
    .A2(net336));
 sg13g2_a21oi_1 _2003_ (.A1(net70),
    .A2(net336),
    .Y(_0037_),
    .B1(_0107_));
 sg13g2_a21oi_1 _2004_ (.A1(net385),
    .A2(_0655_),
    .Y(_0108_),
    .B1(net85));
 sg13g2_o21ai_1 _2005_ (.B1(net383),
    .Y(_0109_),
    .A1(_0585_),
    .A2(_0658_));
 sg13g2_nor2_1 _2006_ (.A(_0108_),
    .B(_0109_),
    .Y(_0038_));
 sg13g2_a21oi_1 _2007_ (.A1(net385),
    .A2(_0657_),
    .Y(_0110_),
    .B1(net74));
 sg13g2_nor2_1 _2008_ (.A(_0670_),
    .B(_0110_),
    .Y(_0039_));
 sg13g2_a21oi_1 _2009_ (.A1(net395),
    .A2(_0602_),
    .Y(_0111_),
    .B1(net81));
 sg13g2_and3_2 _2010_ (.X(_0112_),
    .A(net81),
    .B(net395),
    .C(_0602_));
 sg13g2_nor3_1 _2011_ (.A(_0670_),
    .B(_0111_),
    .C(_0112_),
    .Y(_0040_));
 sg13g2_xnor2_1 _2012_ (.Y(_0113_),
    .A(net90),
    .B(_0112_));
 sg13g2_nor2_1 _2013_ (.A(_0670_),
    .B(_0113_),
    .Y(_0041_));
 sg13g2_a21oi_1 _2014_ (.A1(\u8.rbop[1] ),
    .A2(_0112_),
    .Y(_0114_),
    .B1(net72));
 sg13g2_nor2_1 _2015_ (.A(_0670_),
    .B(net73),
    .Y(_0042_));
 sg13g2_nor4_1 _2016_ (.A(net301),
    .B(net385),
    .C(_0646_),
    .D(_0651_),
    .Y(_0115_));
 sg13g2_o21ai_1 _2017_ (.B1(net383),
    .Y(_0116_),
    .A1(net102),
    .A2(_0115_));
 sg13g2_and2_1 _2018_ (.A(net102),
    .B(_0115_),
    .X(_0117_));
 sg13g2_nor2_1 _2019_ (.A(_0116_),
    .B(_0117_),
    .Y(_0043_));
 sg13g2_o21ai_1 _2020_ (.B1(net383),
    .Y(_0118_),
    .A1(net77),
    .A2(_0117_));
 sg13g2_a21oi_1 _2021_ (.A1(net77),
    .A2(_0117_),
    .Y(_0044_),
    .B1(_0118_));
 sg13g2_a21oi_1 _2022_ (.A1(net77),
    .A2(_0117_),
    .Y(_0119_),
    .B1(net79));
 sg13g2_nor2_1 _2023_ (.A(_0670_),
    .B(net80),
    .Y(_0045_));
 sg13g2_nand2_1 _2024_ (.Y(_0120_),
    .A(net364),
    .B(net305));
 sg13g2_o21ai_1 _2025_ (.B1(_0120_),
    .Y(_0121_),
    .A1(net353),
    .A2(_0576_));
 sg13g2_o21ai_1 _2026_ (.B1(_0458_),
    .Y(_0122_),
    .A1(_0478_),
    .A2(_0121_));
 sg13g2_a22oi_1 _2027_ (.Y(_0123_),
    .B1(net8),
    .B2(_0939_),
    .A2(net413),
    .A1(\u8.ls[8] ));
 sg13g2_nor2_1 _2028_ (.A(_0472_),
    .B(_0123_),
    .Y(_0124_));
 sg13g2_a21oi_1 _2029_ (.A1(net360),
    .A2(net317),
    .Y(_0125_),
    .B1(net325));
 sg13g2_o21ai_1 _2030_ (.B1(_0122_),
    .Y(_0126_),
    .A1(_0451_),
    .A2(_0125_));
 sg13g2_nor3_1 _2031_ (.A(_0937_),
    .B(_0124_),
    .C(_0126_),
    .Y(_0127_));
 sg13g2_o21ai_1 _2032_ (.B1(net417),
    .Y(_0128_),
    .A1(net348),
    .A2(net290));
 sg13g2_nor2_1 _2033_ (.A(_0127_),
    .B(_0128_),
    .Y(_0046_));
 sg13g2_xor2_1 _2034_ (.B(net352),
    .A(net349),
    .X(_0129_));
 sg13g2_a22oi_1 _2035_ (.Y(_0130_),
    .B1(_0575_),
    .B2(_0129_),
    .A2(net304),
    .A1(\u8.ls[9] ));
 sg13g2_nor3_1 _2036_ (.A(net314),
    .B(_0459_),
    .C(_0130_),
    .Y(_0131_));
 sg13g2_nand3_1 _2037_ (.B(_0433_),
    .C(net317),
    .A(net358),
    .Y(_0132_));
 sg13g2_a21oi_1 _2038_ (.A1(net334),
    .A2(_0132_),
    .Y(_0133_),
    .B1(_0451_));
 sg13g2_nor2_1 _2039_ (.A(net413),
    .B(_0930_),
    .Y(_0134_));
 sg13g2_or2_1 _2040_ (.X(_0135_),
    .B(_0134_),
    .A(_0472_));
 sg13g2_nor3_1 _2041_ (.A(_0488_),
    .B(_0686_),
    .C(_0135_),
    .Y(_0136_));
 sg13g2_nor4_1 _2042_ (.A(_0937_),
    .B(_0131_),
    .C(_0133_),
    .D(_0136_),
    .Y(_0137_));
 sg13g2_o21ai_1 _2043_ (.B1(net418),
    .Y(_0138_),
    .A1(net100),
    .A2(net290));
 sg13g2_nor2_1 _2044_ (.A(_0137_),
    .B(_0138_),
    .Y(_0047_));
 sg13g2_xnor2_1 _2045_ (.Y(_0139_),
    .A(_0194_),
    .B(_0228_));
 sg13g2_nor2_1 _2046_ (.A(net314),
    .B(_0139_),
    .Y(_0140_));
 sg13g2_a22oi_1 _2047_ (.Y(_0141_),
    .B1(_0575_),
    .B2(_0140_),
    .A2(net305),
    .A1(net360));
 sg13g2_and3_1 _2048_ (.X(_0142_),
    .A(net335),
    .B(_0433_),
    .C(net316));
 sg13g2_nand2_1 _2049_ (.Y(_0143_),
    .A(net103),
    .B(_0142_));
 sg13g2_a221oi_1 _2050_ (.B2(net310),
    .C1(net386),
    .B1(_0143_),
    .A1(net294),
    .Y(_0144_),
    .A2(_0141_));
 sg13g2_nor3_1 _2051_ (.A(_0498_),
    .B(_0625_),
    .C(_0135_),
    .Y(_0145_));
 sg13g2_nor3_1 _2052_ (.A(_0937_),
    .B(_0144_),
    .C(_0145_),
    .Y(_0146_));
 sg13g2_o21ai_1 _2053_ (.B1(net417),
    .Y(_0147_),
    .A1(net345),
    .A2(net290));
 sg13g2_nor2_1 _2054_ (.A(_0146_),
    .B(_0147_),
    .Y(_0048_));
 sg13g2_xnor2_1 _2055_ (.Y(_0148_),
    .A(_0193_),
    .B(_0317_));
 sg13g2_nor3_1 _2056_ (.A(net314),
    .B(_0572_),
    .C(_0148_),
    .Y(_0149_));
 sg13g2_a21oi_1 _2057_ (.A1(net358),
    .A2(net304),
    .Y(_0150_),
    .B1(_0149_));
 sg13g2_a21o_1 _2058_ (.A2(_0142_),
    .A1(net355),
    .B1(_1011_),
    .X(_0151_));
 sg13g2_a21oi_1 _2059_ (.A1(net294),
    .A2(_0150_),
    .Y(_0152_),
    .B1(net386));
 sg13g2_nor3_1 _2060_ (.A(_0512_),
    .B(_0691_),
    .C(_0135_),
    .Y(_0153_));
 sg13g2_a21oi_1 _2061_ (.A1(_0151_),
    .A2(_0152_),
    .Y(_0154_),
    .B1(_0153_));
 sg13g2_o21ai_1 _2062_ (.B1(net417),
    .Y(_0155_),
    .A1(net344),
    .A2(net290));
 sg13g2_a21oi_1 _2063_ (.A1(net290),
    .A2(_0154_),
    .Y(_0049_),
    .B1(_0155_));
 sg13g2_nor4_1 _2064_ (.A(_0193_),
    .B(_0317_),
    .C(net314),
    .D(_0572_),
    .Y(_0156_));
 sg13g2_a21oi_1 _2065_ (.A1(net356),
    .A2(net304),
    .Y(_0157_),
    .B1(_0156_));
 sg13g2_nand2_1 _2066_ (.Y(_0158_),
    .A(net352),
    .B(_0142_));
 sg13g2_a221oi_1 _2067_ (.B2(net310),
    .C1(net386),
    .B1(_0158_),
    .A1(net294),
    .Y(_0159_),
    .A2(_0157_));
 sg13g2_nor2b_1 _2068_ (.A(_0524_),
    .B_N(_0739_),
    .Y(_0160_));
 sg13g2_o21ai_1 _2069_ (.B1(net290),
    .Y(_0161_),
    .A1(_0135_),
    .A2(_0160_));
 sg13g2_o21ai_1 _2070_ (.B1(net417),
    .Y(_0162_),
    .A1(_0159_),
    .A2(_0161_));
 sg13g2_a21oi_1 _2071_ (.A1(_0190_),
    .A2(_0937_),
    .Y(_0050_),
    .B1(_0162_));
 sg13g2_nand3_1 _2072_ (.B(_0433_),
    .C(net316),
    .A(net350),
    .Y(_0163_));
 sg13g2_a21oi_1 _2073_ (.A1(net335),
    .A2(_0163_),
    .Y(_0164_),
    .B1(_0451_));
 sg13g2_nand2_1 _2074_ (.Y(_0165_),
    .A(net13),
    .B(_0939_));
 sg13g2_a21oi_1 _2075_ (.A1(_0856_),
    .A2(_0165_),
    .Y(_0166_),
    .B1(_0472_));
 sg13g2_nor3_1 _2076_ (.A(_0200_),
    .B(_0459_),
    .C(_0465_),
    .Y(_0167_));
 sg13g2_nor4_1 _2077_ (.A(_0937_),
    .B(_0164_),
    .C(_0166_),
    .D(_0167_),
    .Y(_0168_));
 sg13g2_o21ai_1 _2078_ (.B1(net418),
    .Y(_0169_),
    .A1(net341),
    .A2(_0936_));
 sg13g2_nor2_1 _2079_ (.A(_0168_),
    .B(_0169_),
    .Y(_0051_));
 sg13g2_a21o_1 _2080_ (.A2(net318),
    .A1(net308),
    .B1(net311),
    .X(_0170_));
 sg13g2_a221oi_1 _2081_ (.B2(net347),
    .C1(_0434_),
    .B1(_0170_),
    .A1(_0436_),
    .Y(_0171_),
    .A2(_0803_));
 sg13g2_o21ai_1 _2082_ (.B1(net310),
    .Y(_0172_),
    .A1(net324),
    .A2(_0171_));
 sg13g2_nand2_1 _2083_ (.Y(_0173_),
    .A(net352),
    .B(net304));
 sg13g2_a21oi_1 _2084_ (.A1(net294),
    .A2(_0173_),
    .Y(_0174_),
    .B1(net386));
 sg13g2_nand2b_1 _2085_ (.Y(_0175_),
    .B(_0817_),
    .A_N(_0539_));
 sg13g2_nor2_1 _2086_ (.A(_0135_),
    .B(_0175_),
    .Y(_0176_));
 sg13g2_a21oi_1 _2087_ (.A1(_0172_),
    .A2(_0174_),
    .Y(_0177_),
    .B1(_0176_));
 sg13g2_o21ai_1 _2088_ (.B1(net417),
    .Y(_0178_),
    .A1(net92),
    .A2(net290));
 sg13g2_a21oi_1 _2089_ (.A1(net290),
    .A2(_0177_),
    .Y(_0052_),
    .B1(_0178_));
 sg13g2_nor2b_1 _2090_ (.A(_0547_),
    .B_N(_0847_),
    .Y(_0179_));
 sg13g2_nand2_1 _2091_ (.Y(_0180_),
    .A(\u8.rc[17] ),
    .B(_0424_));
 sg13g2_nand2_1 _2092_ (.Y(_0181_),
    .A(\u8.rc[17] ),
    .B(net316));
 sg13g2_a221oi_1 _2093_ (.B2(net307),
    .C1(net324),
    .B1(_0181_),
    .A1(_0439_),
    .Y(_0182_),
    .A2(_0180_));
 sg13g2_nand2_1 _2094_ (.Y(_0183_),
    .A(net349),
    .B(net304));
 sg13g2_a21oi_1 _2095_ (.A1(net294),
    .A2(_0183_),
    .Y(_0184_),
    .B1(net386));
 sg13g2_o21ai_1 _2096_ (.B1(_0184_),
    .Y(_0185_),
    .A1(_1011_),
    .A2(_0182_));
 sg13g2_o21ai_1 _2097_ (.B1(_0185_),
    .Y(_0186_),
    .A1(_0135_),
    .A2(_0179_));
 sg13g2_o21ai_1 _2098_ (.B1(net417),
    .Y(_0187_),
    .A1(_0937_),
    .A2(_0186_));
 sg13g2_a21oi_1 _2099_ (.A1(_0188_),
    .A2(_0937_),
    .Y(_0053_),
    .B1(_0187_));
 sg13g2_dfrbpq_2 _2100_ (.RESET_B(net46),
    .D(net99),
    .Q(\u8.rc[24] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2101_ (.RESET_B(net35),
    .D(_0001_),
    .Q(\u8.rc[25] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2102_ (.RESET_B(net33),
    .D(_0002_),
    .Q(\u8.rc[26] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _2103_ (.RESET_B(net31),
    .D(_0003_),
    .Q(\u8.rc[27] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _2104_ (.RESET_B(net29),
    .D(_0004_),
    .Q(\u8.rc[28] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2105_ (.RESET_B(net27),
    .D(_0005_),
    .Q(\u8.rc[29] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _2106_ (.RESET_B(net25),
    .D(_0006_),
    .Q(\u8.rc[30] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _2107_ (.RESET_B(net23),
    .D(_0007_),
    .Q(\u8.rc[31] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _2108_ (.RESET_B(net21),
    .D(_0008_),
    .Q(retry),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _2109_ (.RESET_B(net19),
    .D(_0009_),
    .Q(uio_out[0]),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2110_ (.RESET_B(net17),
    .D(_0010_),
    .Q(uio_out[1]),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2111_ (.RESET_B(net69),
    .D(_0011_),
    .Q(uio_out[2]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _2112_ (.RESET_B(net67),
    .D(_0012_),
    .Q(uio_out[3]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _2113_ (.RESET_B(net65),
    .D(_0013_),
    .Q(uio_out[4]),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2114_ (.RESET_B(net63),
    .D(_0014_),
    .Q(uio_out[5]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _2115_ (.RESET_B(net61),
    .D(_0015_),
    .Q(uio_out[6]),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _2116_ (.RESET_B(net59),
    .D(_0016_),
    .Q(uio_out[7]),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _2117_ (.RESET_B(net57),
    .D(_0017_),
    .Q(\u8.empty ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _2118_ (.RESET_B(net55),
    .D(_0018_),
    .Q(\u8.ls[0] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _2119_ (.RESET_B(net53),
    .D(_0019_),
    .Q(\u8.ls[1] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _2120_ (.RESET_B(net51),
    .D(_0020_),
    .Q(\u8.ls[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _2121_ (.RESET_B(net49),
    .D(_0021_),
    .Q(\u8.ls[3] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _2122_ (.RESET_B(net47),
    .D(_0022_),
    .Q(\u8.ls[4] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _2123_ (.RESET_B(net45),
    .D(_0023_),
    .Q(\u8.ls[5] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _2124_ (.RESET_B(net43),
    .D(_0024_),
    .Q(\u8.ls[6] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _2125_ (.RESET_B(net41),
    .D(_0025_),
    .Q(\u8.ls[7] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _2126_ (.RESET_B(net39),
    .D(_0026_),
    .Q(\u8.ls[8] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _2127_ (.RESET_B(net37),
    .D(_0027_),
    .Q(\u8.ls[9] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _2128_ (.RESET_B(net34),
    .D(net118),
    .Q(\u8.hs[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _2129_ (.RESET_B(net30),
    .D(_0029_),
    .Q(\u8.hs[1] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _2130_ (.RESET_B(net26),
    .D(_0030_),
    .Q(\u8.hs[2] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _2131_ (.RESET_B(net22),
    .D(_0031_),
    .Q(\u8.hs[3] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _2132_ (.RESET_B(net18),
    .D(_0032_),
    .Q(\u8.hs[4] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _2133_ (.RESET_B(net68),
    .D(_0033_),
    .Q(\u8.hs[5] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _2134_ (.RESET_B(net64),
    .D(_0034_),
    .Q(\u8.rcip[0] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _2135_ (.RESET_B(net60),
    .D(net83),
    .Q(\u8.rcip[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _2136_ (.RESET_B(net56),
    .D(_0036_),
    .Q(\u8.rcip[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _2137_ (.RESET_B(net52),
    .D(net71),
    .Q(\u8.rcop[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2138_ (.RESET_B(net48),
    .D(_0038_),
    .Q(\u8.rcop[1] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2139_ (.RESET_B(net44),
    .D(_0039_),
    .Q(\u8.rcop[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2140_ (.RESET_B(net40),
    .D(_0040_),
    .Q(\u8.rbop[0] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_2 _2141_ (.RESET_B(net36),
    .D(_0041_),
    .Q(\u8.rbop[1] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _2142_ (.RESET_B(net28),
    .D(_0042_),
    .Q(\u8.rbop[2] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _2143_ (.RESET_B(net20),
    .D(_0043_),
    .Q(\u8.ruop[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _2144_ (.RESET_B(net66),
    .D(net78),
    .Q(\u8.ruop[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _2145_ (.RESET_B(net58),
    .D(_0045_),
    .Q(\u8.ruop[2] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _2146_ (.RESET_B(net50),
    .D(net111),
    .Q(\u8.rc[16] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2147_ (.RESET_B(net42),
    .D(_0047_),
    .Q(\u8.rc[17] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2148_ (.RESET_B(net32),
    .D(_0048_),
    .Q(\u8.rc[18] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _2149_ (.RESET_B(net16),
    .D(_0049_),
    .Q(\u8.rc[19] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _2150_ (.RESET_B(net54),
    .D(_0050_),
    .Q(\u8.rc[20] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _2151_ (.RESET_B(net38),
    .D(_0051_),
    .Q(\u8.rc[21] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _2152_ (.RESET_B(net62),
    .D(_0052_),
    .Q(\u8.rc[22] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_1 _2153_ (.RESET_B(net24),
    .D(_0053_),
    .Q(\u8.rc[23] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_tiehi _2110__17 (.L_HI(net17));
 sg13g2_tiehi _2132__18 (.L_HI(net18));
 sg13g2_tiehi _2109__19 (.L_HI(net19));
 sg13g2_tiehi _2143__20 (.L_HI(net20));
 sg13g2_tiehi _2108__21 (.L_HI(net21));
 sg13g2_tiehi _2131__22 (.L_HI(net22));
 sg13g2_tiehi _2107__23 (.L_HI(net23));
 sg13g2_tiehi _2153__24 (.L_HI(net24));
 sg13g2_tiehi _2106__25 (.L_HI(net25));
 sg13g2_tiehi _2130__26 (.L_HI(net26));
 sg13g2_tiehi _2105__27 (.L_HI(net27));
 sg13g2_tiehi _2142__28 (.L_HI(net28));
 sg13g2_tiehi _2104__29 (.L_HI(net29));
 sg13g2_tiehi _2129__30 (.L_HI(net30));
 sg13g2_tiehi _2103__31 (.L_HI(net31));
 sg13g2_tiehi _2148__32 (.L_HI(net32));
 sg13g2_tiehi _2102__33 (.L_HI(net33));
 sg13g2_tiehi _2128__34 (.L_HI(net34));
 sg13g2_tiehi _2101__35 (.L_HI(net35));
 sg13g2_tiehi _2141__36 (.L_HI(net36));
 sg13g2_tiehi _2127__37 (.L_HI(net37));
 sg13g2_tiehi _2151__38 (.L_HI(net38));
 sg13g2_tiehi _2126__39 (.L_HI(net39));
 sg13g2_tiehi _2140__40 (.L_HI(net40));
 sg13g2_tiehi _2125__41 (.L_HI(net41));
 sg13g2_tiehi _2147__42 (.L_HI(net42));
 sg13g2_tiehi _2124__43 (.L_HI(net43));
 sg13g2_tiehi _2139__44 (.L_HI(net44));
 sg13g2_tiehi _2123__45 (.L_HI(net45));
 sg13g2_tiehi _2100__46 (.L_HI(net46));
 sg13g2_tiehi _2122__47 (.L_HI(net47));
 sg13g2_tiehi _2138__48 (.L_HI(net48));
 sg13g2_tiehi _2121__49 (.L_HI(net49));
 sg13g2_tiehi _2146__50 (.L_HI(net50));
 sg13g2_tiehi _2120__51 (.L_HI(net51));
 sg13g2_tiehi _2137__52 (.L_HI(net52));
 sg13g2_tiehi _2119__53 (.L_HI(net53));
 sg13g2_tiehi _2150__54 (.L_HI(net54));
 sg13g2_tiehi _2118__55 (.L_HI(net55));
 sg13g2_tiehi _2136__56 (.L_HI(net56));
 sg13g2_tiehi _2117__57 (.L_HI(net57));
 sg13g2_tiehi _2145__58 (.L_HI(net58));
 sg13g2_tiehi _2116__59 (.L_HI(net59));
 sg13g2_tiehi _2135__60 (.L_HI(net60));
 sg13g2_tiehi _2115__61 (.L_HI(net61));
 sg13g2_tiehi _2152__62 (.L_HI(net62));
 sg13g2_tiehi _2114__63 (.L_HI(net63));
 sg13g2_tiehi _2134__64 (.L_HI(net64));
 sg13g2_tiehi _2113__65 (.L_HI(net65));
 sg13g2_tiehi _2144__66 (.L_HI(net66));
 sg13g2_tiehi _2112__67 (.L_HI(net67));
 sg13g2_tiehi _2133__68 (.L_HI(net68));
 sg13g2_tiehi _2111__69 (.L_HI(net69));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _2208_ (.A(net397),
    .X(uio_oe[0]));
 sg13g2_buf_1 _2209_ (.A(net397),
    .X(uio_oe[1]));
 sg13g2_buf_1 _2210_ (.A(net397),
    .X(uio_oe[2]));
 sg13g2_buf_1 _2211_ (.A(net396),
    .X(uio_oe[3]));
 sg13g2_buf_1 _2212_ (.A(net396),
    .X(uio_oe[4]));
 sg13g2_buf_1 _2213_ (.A(net396),
    .X(uio_oe[5]));
 sg13g2_buf_1 _2214_ (.A(net396),
    .X(uio_oe[6]));
 sg13g2_buf_1 _2215_ (.A(net397),
    .X(uio_oe[7]));
 sg13g2_buf_8 fanout285 (.A(net287),
    .X(net285));
 sg13g2_buf_1 fanout286 (.A(net287),
    .X(net286));
 sg13g2_buf_8 fanout287 (.A(_0940_),
    .X(net287));
 sg13g2_buf_8 fanout288 (.A(net289),
    .X(net288));
 sg13g2_buf_8 fanout289 (.A(_0940_),
    .X(net289));
 sg13g2_buf_8 fanout290 (.A(_0936_),
    .X(net290));
 sg13g2_buf_8 fanout291 (.A(_0469_),
    .X(net291));
 sg13g2_buf_8 fanout292 (.A(_0947_),
    .X(net292));
 sg13g2_buf_8 fanout293 (.A(_0946_),
    .X(net293));
 sg13g2_buf_8 fanout294 (.A(net296),
    .X(net294));
 sg13g2_buf_8 fanout295 (.A(net296),
    .X(net295));
 sg13g2_buf_2 fanout296 (.A(_0944_),
    .X(net296));
 sg13g2_buf_2 fanout297 (.A(_0586_),
    .X(net297));
 sg13g2_buf_1 fanout298 (.A(_0586_),
    .X(net298));
 sg13g2_buf_8 fanout299 (.A(_0415_),
    .X(net299));
 sg13g2_buf_8 fanout300 (.A(_0415_),
    .X(net300));
 sg13g2_buf_8 fanout301 (.A(_0390_),
    .X(net301));
 sg13g2_buf_8 fanout302 (.A(_0573_),
    .X(net302));
 sg13g2_buf_8 fanout303 (.A(_0465_),
    .X(net303));
 sg13g2_buf_8 fanout304 (.A(net305),
    .X(net304));
 sg13g2_buf_8 fanout305 (.A(net306),
    .X(net305));
 sg13g2_buf_8 fanout306 (.A(_0464_),
    .X(net306));
 sg13g2_buf_8 fanout307 (.A(net308),
    .X(net307));
 sg13g2_buf_8 fanout308 (.A(_0430_),
    .X(net308));
 sg13g2_buf_8 fanout309 (.A(_0477_),
    .X(net309));
 sg13g2_buf_8 fanout310 (.A(_1010_),
    .X(net310));
 sg13g2_buf_8 fanout311 (.A(_0424_),
    .X(net311));
 sg13g2_buf_8 fanout312 (.A(_0412_),
    .X(net312));
 sg13g2_buf_8 fanout313 (.A(_0384_),
    .X(net313));
 sg13g2_buf_1 fanout314 (.A(_0384_),
    .X(net314));
 sg13g2_buf_8 fanout315 (.A(_0452_),
    .X(net315));
 sg13g2_buf_8 fanout316 (.A(net318),
    .X(net316));
 sg13g2_buf_1 fanout317 (.A(net318),
    .X(net317));
 sg13g2_buf_8 fanout318 (.A(_0442_),
    .X(net318));
 sg13g2_buf_8 fanout319 (.A(_0396_),
    .X(net319));
 sg13g2_buf_8 fanout320 (.A(_0379_),
    .X(net320));
 sg13g2_buf_8 fanout321 (.A(_0993_),
    .X(net321));
 sg13g2_buf_8 fanout322 (.A(_0635_),
    .X(net322));
 sg13g2_buf_8 fanout323 (.A(_0473_),
    .X(net323));
 sg13g2_buf_8 fanout324 (.A(net325),
    .X(net324));
 sg13g2_buf_8 fanout325 (.A(_0395_),
    .X(net325));
 sg13g2_buf_8 fanout326 (.A(_0660_),
    .X(net326));
 sg13g2_buf_8 fanout327 (.A(net328),
    .X(net327));
 sg13g2_buf_8 fanout328 (.A(_0618_),
    .X(net328));
 sg13g2_buf_8 fanout329 (.A(_0616_),
    .X(net329));
 sg13g2_buf_8 fanout330 (.A(_0615_),
    .X(net330));
 sg13g2_buf_1 fanout331 (.A(_0615_),
    .X(net331));
 sg13g2_buf_8 fanout332 (.A(net333),
    .X(net332));
 sg13g2_buf_8 fanout333 (.A(_0615_),
    .X(net333));
 sg13g2_buf_8 fanout334 (.A(net335),
    .X(net334));
 sg13g2_buf_8 fanout335 (.A(_0394_),
    .X(net335));
 sg13g2_buf_8 fanout336 (.A(_0665_),
    .X(net336));
 sg13g2_buf_8 fanout337 (.A(_0211_),
    .X(net337));
 sg13g2_buf_8 fanout338 (.A(net113),
    .X(net338));
 sg13g2_buf_8 fanout339 (.A(\u8.rc[22] ),
    .X(net339));
 sg13g2_buf_8 fanout340 (.A(\u8.rc[21] ),
    .X(net340));
 sg13g2_buf_8 fanout341 (.A(net116),
    .X(net341));
 sg13g2_buf_8 fanout342 (.A(net120),
    .X(net342));
 sg13g2_buf_8 fanout343 (.A(\u8.rc[19] ),
    .X(net343));
 sg13g2_buf_1 fanout344 (.A(net124),
    .X(net344));
 sg13g2_buf_8 fanout345 (.A(net130),
    .X(net345));
 sg13g2_buf_8 fanout346 (.A(\u8.rc[17] ),
    .X(net346));
 sg13g2_buf_8 fanout347 (.A(net348),
    .X(net347));
 sg13g2_buf_8 fanout348 (.A(net110),
    .X(net348));
 sg13g2_buf_8 fanout349 (.A(\u8.hs[5] ),
    .X(net349));
 sg13g2_buf_8 fanout350 (.A(net119),
    .X(net350));
 sg13g2_buf_8 fanout351 (.A(net353),
    .X(net351));
 sg13g2_buf_8 fanout352 (.A(net353),
    .X(net352));
 sg13g2_buf_8 fanout353 (.A(net131),
    .X(net353));
 sg13g2_buf_8 fanout354 (.A(\u8.hs[3] ),
    .X(net354));
 sg13g2_buf_2 fanout355 (.A(net129),
    .X(net355));
 sg13g2_buf_8 fanout356 (.A(\u8.hs[2] ),
    .X(net356));
 sg13g2_buf_8 fanout357 (.A(\u8.hs[1] ),
    .X(net357));
 sg13g2_buf_8 fanout358 (.A(net112),
    .X(net358));
 sg13g2_buf_8 fanout359 (.A(\u8.hs[0] ),
    .X(net359));
 sg13g2_buf_8 fanout360 (.A(net117),
    .X(net360));
 sg13g2_buf_8 fanout361 (.A(net127),
    .X(net361));
 sg13g2_buf_8 fanout362 (.A(\u8.ls[9] ),
    .X(net362));
 sg13g2_buf_8 fanout363 (.A(net364),
    .X(net363));
 sg13g2_buf_8 fanout364 (.A(net122),
    .X(net364));
 sg13g2_buf_8 fanout365 (.A(net367),
    .X(net365));
 sg13g2_buf_1 fanout366 (.A(net367),
    .X(net366));
 sg13g2_buf_8 fanout367 (.A(net107),
    .X(net367));
 sg13g2_buf_8 fanout368 (.A(net369),
    .X(net368));
 sg13g2_buf_8 fanout369 (.A(net121),
    .X(net369));
 sg13g2_buf_8 fanout370 (.A(\u8.ls[5] ),
    .X(net370));
 sg13g2_buf_8 fanout371 (.A(net114),
    .X(net371));
 sg13g2_buf_1 fanout372 (.A(\u8.ls[4] ),
    .X(net372));
 sg13g2_buf_8 fanout373 (.A(\u8.ls[2] ),
    .X(net373));
 sg13g2_buf_8 fanout374 (.A(net123),
    .X(net374));
 sg13g2_buf_8 fanout375 (.A(net128),
    .X(net375));
 sg13g2_buf_8 fanout376 (.A(net377),
    .X(net376));
 sg13g2_buf_8 fanout377 (.A(\u8.rc[31] ),
    .X(net377));
 sg13g2_buf_8 fanout378 (.A(\u8.rc[30] ),
    .X(net378));
 sg13g2_buf_8 fanout379 (.A(net126),
    .X(net379));
 sg13g2_buf_8 fanout380 (.A(net125),
    .X(net380));
 sg13g2_buf_8 fanout381 (.A(net115),
    .X(net381));
 sg13g2_buf_8 fanout382 (.A(\u8.rc[24] ),
    .X(net382));
 sg13g2_buf_8 fanout383 (.A(_0669_),
    .X(net383));
 sg13g2_buf_1 fanout384 (.A(_0669_),
    .X(net384));
 sg13g2_buf_8 fanout385 (.A(_0584_),
    .X(net385));
 sg13g2_buf_8 fanout386 (.A(_0449_),
    .X(net386));
 sg13g2_buf_1 fanout387 (.A(_0449_),
    .X(net387));
 sg13g2_buf_2 fanout388 (.A(net389),
    .X(net388));
 sg13g2_buf_1 fanout389 (.A(net390),
    .X(net389));
 sg13g2_buf_1 fanout390 (.A(_0449_),
    .X(net390));
 sg13g2_buf_8 fanout391 (.A(net392),
    .X(net391));
 sg13g2_buf_8 fanout392 (.A(_0222_),
    .X(net392));
 sg13g2_buf_8 fanout393 (.A(net394),
    .X(net393));
 sg13g2_buf_8 fanout394 (.A(_0222_),
    .X(net394));
 sg13g2_buf_8 fanout395 (.A(net5),
    .X(net395));
 sg13g2_buf_2 fanout396 (.A(net397),
    .X(net396));
 sg13g2_buf_1 fanout397 (.A(net398),
    .X(net397));
 sg13g2_buf_1 fanout398 (.A(net399),
    .X(net398));
 sg13g2_buf_8 fanout399 (.A(net4),
    .X(net399));
 sg13g2_buf_8 fanout400 (.A(net402),
    .X(net400));
 sg13g2_buf_2 fanout401 (.A(net402),
    .X(net401));
 sg13g2_buf_8 fanout402 (.A(net406),
    .X(net402));
 sg13g2_buf_8 fanout403 (.A(net404),
    .X(net403));
 sg13g2_buf_8 fanout404 (.A(net405),
    .X(net404));
 sg13g2_buf_8 fanout405 (.A(net406),
    .X(net405));
 sg13g2_buf_8 fanout406 (.A(net415),
    .X(net406));
 sg13g2_buf_8 fanout407 (.A(net408),
    .X(net407));
 sg13g2_buf_8 fanout408 (.A(net415),
    .X(net408));
 sg13g2_buf_8 fanout409 (.A(net411),
    .X(net409));
 sg13g2_buf_1 fanout410 (.A(net411),
    .X(net410));
 sg13g2_buf_1 fanout411 (.A(net415),
    .X(net411));
 sg13g2_buf_8 fanout412 (.A(net414),
    .X(net412));
 sg13g2_buf_1 fanout413 (.A(net414),
    .X(net413));
 sg13g2_buf_1 fanout414 (.A(net415),
    .X(net414));
 sg13g2_buf_2 fanout415 (.A(ui_in[3]),
    .X(net415));
 sg13g2_buf_8 fanout416 (.A(net421),
    .X(net416));
 sg13g2_buf_8 fanout417 (.A(net421),
    .X(net417));
 sg13g2_buf_1 fanout418 (.A(net421),
    .X(net418));
 sg13g2_buf_8 fanout419 (.A(net420),
    .X(net419));
 sg13g2_buf_8 fanout420 (.A(net421),
    .X(net420));
 sg13g2_buf_8 fanout421 (.A(rst_n),
    .X(net421));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[6]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(ui_in[7]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[0]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[1]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[2]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[3]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[4]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[5]),
    .X(net13));
 sg13g2_buf_1 input14 (.A(uio_in[6]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[7]),
    .X(net15));
 sg13g2_tiehi _2149__16 (.L_HI(net16));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_inv_1 clkload2 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_4__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_5__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_6__leaf_clk));
 sg13g2_inv_1 clkload6 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\u8.rcop[0] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0037_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold3 (.A(\u8.rbop[2] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0114_),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold5 (.A(\u8.rcop[2] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold6 (.A(\u8.rcip[0] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0102_),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold8 (.A(\u8.ruop[1] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold9 (.A(_0044_),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold10 (.A(\u8.ruop[2] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0119_),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold12 (.A(\u8.rbop[0] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold13 (.A(\u8.rcip[1] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold14 (.A(_0035_),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold15 (.A(\u8.rcip[2] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold16 (.A(\u8.rcop[1] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold17 (.A(uio_out[6]),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold18 (.A(uio_out[1]),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold19 (.A(uio_out[0]),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold20 (.A(uio_out[4]),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold21 (.A(\u8.rbop[1] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold22 (.A(uio_out[7]),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold23 (.A(\u8.rc[22] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold24 (.A(uio_out[5]),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold25 (.A(uio_out[3]),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold26 (.A(uio_out[2]),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold27 (.A(\u8.rc[30] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold28 (.A(retry),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold29 (.A(\u8.rc[24] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold30 (.A(_0000_),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold31 (.A(\u8.rc[17] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold32 (.A(\u8.ls[2] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold33 (.A(\u8.ruop[0] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold34 (.A(\u8.hs[2] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold35 (.A(\u8.ls[5] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold36 (.A(\u8.rc[28] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold37 (.A(\u8.rc[26] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold38 (.A(\u8.ls[7] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold39 (.A(\u8.ls[0] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold40 (.A(\u8.ls[3] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold41 (.A(\u8.rc[16] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0046_),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold43 (.A(\u8.hs[1] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold44 (.A(\u8.rc[23] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold45 (.A(\u8.ls[4] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold46 (.A(\u8.rc[25] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold47 (.A(\u8.rc[21] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold48 (.A(\u8.hs[0] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0028_),
    .X(net118));
 sg13g2_dlygate4sd3_1 hold50 (.A(\u8.hs[5] ),
    .X(net119));
 sg13g2_dlygate4sd3_1 hold51 (.A(\u8.rc[20] ),
    .X(net120));
 sg13g2_dlygate4sd3_1 hold52 (.A(\u8.ls[6] ),
    .X(net121));
 sg13g2_dlygate4sd3_1 hold53 (.A(\u8.ls[8] ),
    .X(net122));
 sg13g2_dlygate4sd3_1 hold54 (.A(\u8.ls[1] ),
    .X(net123));
 sg13g2_dlygate4sd3_1 hold55 (.A(\u8.rc[19] ),
    .X(net124));
 sg13g2_dlygate4sd3_1 hold56 (.A(\u8.rc[27] ),
    .X(net125));
 sg13g2_dlygate4sd3_1 hold57 (.A(\u8.rc[29] ),
    .X(net126));
 sg13g2_dlygate4sd3_1 hold58 (.A(\u8.ls[9] ),
    .X(net127));
 sg13g2_dlygate4sd3_1 hold59 (.A(\u8.empty ),
    .X(net128));
 sg13g2_dlygate4sd3_1 hold60 (.A(\u8.hs[3] ),
    .X(net129));
 sg13g2_dlygate4sd3_1 hold61 (.A(\u8.rc[18] ),
    .X(net130));
 sg13g2_dlygate4sd3_1 hold62 (.A(\u8.hs[4] ),
    .X(net131));
 sg13g2_dlygate4sd3_1 hold63 (.A(\u8.rc[29] ),
    .X(net132));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_fill_2 FILLER_0_406 ();
 sg13g2_fill_1 FILLER_0_408 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_fill_2 FILLER_1_406 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_8 FILLER_2_203 ();
 sg13g2_decap_8 FILLER_2_210 ();
 sg13g2_decap_8 FILLER_2_217 ();
 sg13g2_decap_8 FILLER_2_224 ();
 sg13g2_decap_8 FILLER_2_231 ();
 sg13g2_decap_8 FILLER_2_238 ();
 sg13g2_decap_8 FILLER_2_245 ();
 sg13g2_decap_8 FILLER_2_252 ();
 sg13g2_decap_8 FILLER_2_259 ();
 sg13g2_decap_8 FILLER_2_266 ();
 sg13g2_decap_8 FILLER_2_273 ();
 sg13g2_decap_8 FILLER_2_280 ();
 sg13g2_decap_8 FILLER_2_287 ();
 sg13g2_decap_8 FILLER_2_294 ();
 sg13g2_decap_8 FILLER_2_301 ();
 sg13g2_decap_8 FILLER_2_308 ();
 sg13g2_decap_8 FILLER_2_315 ();
 sg13g2_decap_8 FILLER_2_322 ();
 sg13g2_decap_8 FILLER_2_329 ();
 sg13g2_decap_8 FILLER_2_336 ();
 sg13g2_decap_8 FILLER_2_343 ();
 sg13g2_decap_8 FILLER_2_350 ();
 sg13g2_decap_8 FILLER_2_357 ();
 sg13g2_decap_8 FILLER_2_364 ();
 sg13g2_decap_8 FILLER_2_371 ();
 sg13g2_decap_8 FILLER_2_378 ();
 sg13g2_decap_8 FILLER_2_385 ();
 sg13g2_decap_8 FILLER_2_392 ();
 sg13g2_decap_8 FILLER_2_399 ();
 sg13g2_fill_2 FILLER_2_406 ();
 sg13g2_fill_1 FILLER_2_408 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_fill_2 FILLER_4_406 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_decap_8 FILLER_5_196 ();
 sg13g2_decap_8 FILLER_5_203 ();
 sg13g2_decap_8 FILLER_5_210 ();
 sg13g2_decap_8 FILLER_5_217 ();
 sg13g2_decap_8 FILLER_5_224 ();
 sg13g2_decap_8 FILLER_5_231 ();
 sg13g2_decap_8 FILLER_5_238 ();
 sg13g2_decap_8 FILLER_5_245 ();
 sg13g2_decap_8 FILLER_5_252 ();
 sg13g2_decap_8 FILLER_5_259 ();
 sg13g2_decap_8 FILLER_5_266 ();
 sg13g2_decap_8 FILLER_5_273 ();
 sg13g2_decap_8 FILLER_5_280 ();
 sg13g2_decap_8 FILLER_5_287 ();
 sg13g2_decap_8 FILLER_5_294 ();
 sg13g2_decap_8 FILLER_5_301 ();
 sg13g2_decap_8 FILLER_5_308 ();
 sg13g2_decap_8 FILLER_5_315 ();
 sg13g2_decap_8 FILLER_5_322 ();
 sg13g2_decap_8 FILLER_5_329 ();
 sg13g2_decap_8 FILLER_5_336 ();
 sg13g2_decap_8 FILLER_5_343 ();
 sg13g2_decap_8 FILLER_5_350 ();
 sg13g2_decap_8 FILLER_5_357 ();
 sg13g2_decap_8 FILLER_5_364 ();
 sg13g2_decap_8 FILLER_5_371 ();
 sg13g2_decap_8 FILLER_5_378 ();
 sg13g2_decap_8 FILLER_5_385 ();
 sg13g2_decap_8 FILLER_5_392 ();
 sg13g2_decap_8 FILLER_5_399 ();
 sg13g2_fill_2 FILLER_5_406 ();
 sg13g2_fill_1 FILLER_5_408 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_fill_2 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_fill_2 FILLER_6_189 ();
 sg13g2_fill_1 FILLER_6_191 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_4 FILLER_6_203 ();
 sg13g2_fill_2 FILLER_6_220 ();
 sg13g2_decap_8 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_247 ();
 sg13g2_fill_1 FILLER_6_249 ();
 sg13g2_decap_8 FILLER_6_254 ();
 sg13g2_decap_8 FILLER_6_261 ();
 sg13g2_decap_8 FILLER_6_268 ();
 sg13g2_decap_8 FILLER_6_275 ();
 sg13g2_decap_8 FILLER_6_282 ();
 sg13g2_decap_8 FILLER_6_289 ();
 sg13g2_decap_8 FILLER_6_296 ();
 sg13g2_decap_8 FILLER_6_303 ();
 sg13g2_decap_8 FILLER_6_310 ();
 sg13g2_decap_8 FILLER_6_317 ();
 sg13g2_decap_8 FILLER_6_324 ();
 sg13g2_decap_8 FILLER_6_331 ();
 sg13g2_decap_8 FILLER_6_338 ();
 sg13g2_decap_8 FILLER_6_345 ();
 sg13g2_decap_8 FILLER_6_352 ();
 sg13g2_decap_8 FILLER_6_359 ();
 sg13g2_decap_8 FILLER_6_366 ();
 sg13g2_decap_8 FILLER_6_373 ();
 sg13g2_decap_8 FILLER_6_380 ();
 sg13g2_decap_8 FILLER_6_387 ();
 sg13g2_decap_8 FILLER_6_394 ();
 sg13g2_decap_8 FILLER_6_401 ();
 sg13g2_fill_1 FILLER_6_408 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_fill_1 FILLER_7_186 ();
 sg13g2_decap_4 FILLER_7_214 ();
 sg13g2_fill_1 FILLER_7_218 ();
 sg13g2_fill_1 FILLER_7_275 ();
 sg13g2_fill_1 FILLER_7_280 ();
 sg13g2_decap_8 FILLER_7_290 ();
 sg13g2_decap_8 FILLER_7_297 ();
 sg13g2_decap_8 FILLER_7_304 ();
 sg13g2_decap_8 FILLER_7_311 ();
 sg13g2_decap_8 FILLER_7_318 ();
 sg13g2_decap_8 FILLER_7_325 ();
 sg13g2_decap_8 FILLER_7_332 ();
 sg13g2_decap_8 FILLER_7_339 ();
 sg13g2_decap_8 FILLER_7_346 ();
 sg13g2_decap_8 FILLER_7_353 ();
 sg13g2_decap_8 FILLER_7_360 ();
 sg13g2_decap_8 FILLER_7_367 ();
 sg13g2_decap_8 FILLER_7_374 ();
 sg13g2_decap_8 FILLER_7_381 ();
 sg13g2_decap_8 FILLER_7_388 ();
 sg13g2_decap_8 FILLER_7_395 ();
 sg13g2_decap_8 FILLER_7_402 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_fill_1 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_89 ();
 sg13g2_decap_8 FILLER_8_96 ();
 sg13g2_decap_8 FILLER_8_103 ();
 sg13g2_decap_8 FILLER_8_110 ();
 sg13g2_decap_8 FILLER_8_117 ();
 sg13g2_decap_4 FILLER_8_137 ();
 sg13g2_fill_1 FILLER_8_141 ();
 sg13g2_decap_8 FILLER_8_146 ();
 sg13g2_fill_1 FILLER_8_158 ();
 sg13g2_decap_4 FILLER_8_177 ();
 sg13g2_decap_4 FILLER_8_192 ();
 sg13g2_decap_4 FILLER_8_209 ();
 sg13g2_decap_4 FILLER_8_226 ();
 sg13g2_decap_8 FILLER_8_299 ();
 sg13g2_decap_8 FILLER_8_306 ();
 sg13g2_decap_8 FILLER_8_313 ();
 sg13g2_decap_8 FILLER_8_320 ();
 sg13g2_decap_8 FILLER_8_327 ();
 sg13g2_decap_8 FILLER_8_334 ();
 sg13g2_decap_8 FILLER_8_341 ();
 sg13g2_decap_8 FILLER_8_348 ();
 sg13g2_decap_8 FILLER_8_355 ();
 sg13g2_decap_8 FILLER_8_362 ();
 sg13g2_decap_8 FILLER_8_369 ();
 sg13g2_decap_8 FILLER_8_376 ();
 sg13g2_decap_8 FILLER_8_383 ();
 sg13g2_decap_8 FILLER_8_390 ();
 sg13g2_decap_8 FILLER_8_397 ();
 sg13g2_decap_4 FILLER_8_404 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_fill_2 FILLER_9_77 ();
 sg13g2_fill_1 FILLER_9_79 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_fill_2 FILLER_9_142 ();
 sg13g2_fill_2 FILLER_9_148 ();
 sg13g2_fill_1 FILLER_9_173 ();
 sg13g2_fill_2 FILLER_9_191 ();
 sg13g2_fill_1 FILLER_9_193 ();
 sg13g2_decap_8 FILLER_9_199 ();
 sg13g2_fill_1 FILLER_9_206 ();
 sg13g2_fill_2 FILLER_9_213 ();
 sg13g2_fill_2 FILLER_9_225 ();
 sg13g2_fill_1 FILLER_9_243 ();
 sg13g2_decap_8 FILLER_9_275 ();
 sg13g2_fill_2 FILLER_9_282 ();
 sg13g2_fill_1 FILLER_9_284 ();
 sg13g2_decap_8 FILLER_9_320 ();
 sg13g2_decap_8 FILLER_9_327 ();
 sg13g2_decap_8 FILLER_9_334 ();
 sg13g2_decap_8 FILLER_9_341 ();
 sg13g2_decap_8 FILLER_9_348 ();
 sg13g2_decap_8 FILLER_9_355 ();
 sg13g2_decap_8 FILLER_9_362 ();
 sg13g2_decap_8 FILLER_9_369 ();
 sg13g2_decap_8 FILLER_9_376 ();
 sg13g2_decap_8 FILLER_9_383 ();
 sg13g2_decap_8 FILLER_9_390 ();
 sg13g2_decap_8 FILLER_9_397 ();
 sg13g2_decap_4 FILLER_9_404 ();
 sg13g2_fill_1 FILLER_9_408 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_decap_8 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_49 ();
 sg13g2_decap_8 FILLER_10_56 ();
 sg13g2_decap_8 FILLER_10_63 ();
 sg13g2_fill_1 FILLER_10_70 ();
 sg13g2_decap_8 FILLER_10_75 ();
 sg13g2_decap_8 FILLER_10_82 ();
 sg13g2_decap_4 FILLER_10_89 ();
 sg13g2_fill_2 FILLER_10_93 ();
 sg13g2_fill_2 FILLER_10_136 ();
 sg13g2_fill_1 FILLER_10_138 ();
 sg13g2_decap_8 FILLER_10_154 ();
 sg13g2_decap_4 FILLER_10_161 ();
 sg13g2_fill_1 FILLER_10_170 ();
 sg13g2_decap_4 FILLER_10_176 ();
 sg13g2_fill_1 FILLER_10_180 ();
 sg13g2_fill_2 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_196 ();
 sg13g2_fill_2 FILLER_10_205 ();
 sg13g2_fill_1 FILLER_10_207 ();
 sg13g2_fill_2 FILLER_10_221 ();
 sg13g2_fill_1 FILLER_10_223 ();
 sg13g2_fill_1 FILLER_10_229 ();
 sg13g2_fill_1 FILLER_10_247 ();
 sg13g2_fill_1 FILLER_10_263 ();
 sg13g2_fill_2 FILLER_10_282 ();
 sg13g2_fill_1 FILLER_10_284 ();
 sg13g2_fill_1 FILLER_10_336 ();
 sg13g2_decap_8 FILLER_10_341 ();
 sg13g2_decap_8 FILLER_10_348 ();
 sg13g2_decap_8 FILLER_10_355 ();
 sg13g2_decap_8 FILLER_10_362 ();
 sg13g2_decap_8 FILLER_10_369 ();
 sg13g2_decap_8 FILLER_10_376 ();
 sg13g2_decap_8 FILLER_10_383 ();
 sg13g2_decap_8 FILLER_10_390 ();
 sg13g2_decap_8 FILLER_10_397 ();
 sg13g2_decap_4 FILLER_10_404 ();
 sg13g2_fill_1 FILLER_10_408 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_fill_2 FILLER_11_63 ();
 sg13g2_fill_1 FILLER_11_65 ();
 sg13g2_fill_1 FILLER_11_94 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_decap_8 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_137 ();
 sg13g2_fill_1 FILLER_11_139 ();
 sg13g2_decap_8 FILLER_11_159 ();
 sg13g2_fill_2 FILLER_11_166 ();
 sg13g2_fill_1 FILLER_11_180 ();
 sg13g2_decap_4 FILLER_11_206 ();
 sg13g2_fill_1 FILLER_11_210 ();
 sg13g2_fill_1 FILLER_11_220 ();
 sg13g2_fill_2 FILLER_11_226 ();
 sg13g2_fill_2 FILLER_11_239 ();
 sg13g2_fill_1 FILLER_11_241 ();
 sg13g2_fill_2 FILLER_11_261 ();
 sg13g2_fill_1 FILLER_11_263 ();
 sg13g2_decap_4 FILLER_11_280 ();
 sg13g2_fill_2 FILLER_11_284 ();
 sg13g2_fill_2 FILLER_11_299 ();
 sg13g2_decap_8 FILLER_11_363 ();
 sg13g2_decap_8 FILLER_11_370 ();
 sg13g2_decap_8 FILLER_11_377 ();
 sg13g2_decap_8 FILLER_11_384 ();
 sg13g2_decap_8 FILLER_11_391 ();
 sg13g2_decap_8 FILLER_11_398 ();
 sg13g2_decap_4 FILLER_11_405 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_decap_8 FILLER_12_28 ();
 sg13g2_decap_8 FILLER_12_35 ();
 sg13g2_decap_8 FILLER_12_42 ();
 sg13g2_decap_8 FILLER_12_49 ();
 sg13g2_decap_4 FILLER_12_84 ();
 sg13g2_fill_2 FILLER_12_88 ();
 sg13g2_decap_4 FILLER_12_95 ();
 sg13g2_fill_2 FILLER_12_115 ();
 sg13g2_decap_8 FILLER_12_128 ();
 sg13g2_fill_2 FILLER_12_135 ();
 sg13g2_fill_1 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_161 ();
 sg13g2_fill_2 FILLER_12_168 ();
 sg13g2_fill_1 FILLER_12_170 ();
 sg13g2_decap_8 FILLER_12_180 ();
 sg13g2_fill_2 FILLER_12_187 ();
 sg13g2_fill_1 FILLER_12_189 ();
 sg13g2_decap_8 FILLER_12_204 ();
 sg13g2_decap_8 FILLER_12_211 ();
 sg13g2_fill_1 FILLER_12_218 ();
 sg13g2_fill_1 FILLER_12_227 ();
 sg13g2_decap_8 FILLER_12_237 ();
 sg13g2_decap_8 FILLER_12_244 ();
 sg13g2_decap_4 FILLER_12_264 ();
 sg13g2_fill_1 FILLER_12_268 ();
 sg13g2_decap_4 FILLER_12_282 ();
 sg13g2_fill_1 FILLER_12_286 ();
 sg13g2_fill_2 FILLER_12_327 ();
 sg13g2_fill_2 FILLER_12_334 ();
 sg13g2_decap_8 FILLER_12_377 ();
 sg13g2_decap_8 FILLER_12_384 ();
 sg13g2_decap_8 FILLER_12_391 ();
 sg13g2_decap_8 FILLER_12_398 ();
 sg13g2_decap_4 FILLER_12_405 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_fill_1 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_66 ();
 sg13g2_decap_4 FILLER_13_73 ();
 sg13g2_fill_2 FILLER_13_99 ();
 sg13g2_fill_1 FILLER_13_101 ();
 sg13g2_fill_2 FILLER_13_117 ();
 sg13g2_decap_8 FILLER_13_132 ();
 sg13g2_decap_4 FILLER_13_158 ();
 sg13g2_fill_2 FILLER_13_162 ();
 sg13g2_decap_8 FILLER_13_184 ();
 sg13g2_decap_4 FILLER_13_191 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_2 FILLER_13_241 ();
 sg13g2_fill_1 FILLER_13_243 ();
 sg13g2_fill_2 FILLER_13_250 ();
 sg13g2_fill_1 FILLER_13_252 ();
 sg13g2_fill_2 FILLER_13_284 ();
 sg13g2_fill_1 FILLER_13_292 ();
 sg13g2_fill_1 FILLER_13_302 ();
 sg13g2_fill_2 FILLER_13_373 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_fill_2 FILLER_13_406 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_4 FILLER_14_42 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_fill_1 FILLER_14_87 ();
 sg13g2_decap_8 FILLER_14_132 ();
 sg13g2_fill_2 FILLER_14_139 ();
 sg13g2_decap_8 FILLER_14_166 ();
 sg13g2_decap_8 FILLER_14_173 ();
 sg13g2_fill_2 FILLER_14_180 ();
 sg13g2_fill_1 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_218 ();
 sg13g2_decap_8 FILLER_14_225 ();
 sg13g2_fill_2 FILLER_14_232 ();
 sg13g2_decap_8 FILLER_14_239 ();
 sg13g2_decap_8 FILLER_14_246 ();
 sg13g2_fill_2 FILLER_14_257 ();
 sg13g2_fill_1 FILLER_14_259 ();
 sg13g2_decap_4 FILLER_14_264 ();
 sg13g2_fill_2 FILLER_14_347 ();
 sg13g2_fill_1 FILLER_14_349 ();
 sg13g2_decap_4 FILLER_14_405 ();
 sg13g2_decap_4 FILLER_15_0 ();
 sg13g2_fill_2 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_34 ();
 sg13g2_fill_2 FILLER_15_41 ();
 sg13g2_decap_8 FILLER_15_50 ();
 sg13g2_decap_8 FILLER_15_57 ();
 sg13g2_fill_1 FILLER_15_64 ();
 sg13g2_fill_1 FILLER_15_81 ();
 sg13g2_fill_2 FILLER_15_99 ();
 sg13g2_fill_1 FILLER_15_106 ();
 sg13g2_fill_1 FILLER_15_113 ();
 sg13g2_decap_8 FILLER_15_147 ();
 sg13g2_decap_4 FILLER_15_154 ();
 sg13g2_fill_1 FILLER_15_158 ();
 sg13g2_fill_1 FILLER_15_169 ();
 sg13g2_fill_2 FILLER_15_178 ();
 sg13g2_decap_4 FILLER_15_185 ();
 sg13g2_fill_1 FILLER_15_206 ();
 sg13g2_decap_4 FILLER_15_216 ();
 sg13g2_decap_4 FILLER_15_232 ();
 sg13g2_fill_2 FILLER_15_236 ();
 sg13g2_decap_8 FILLER_15_253 ();
 sg13g2_decap_4 FILLER_15_260 ();
 sg13g2_fill_2 FILLER_15_264 ();
 sg13g2_fill_2 FILLER_15_281 ();
 sg13g2_fill_1 FILLER_15_283 ();
 sg13g2_fill_2 FILLER_15_315 ();
 sg13g2_fill_1 FILLER_15_332 ();
 sg13g2_fill_2 FILLER_15_375 ();
 sg13g2_fill_1 FILLER_15_377 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_fill_2 FILLER_16_7 ();
 sg13g2_fill_1 FILLER_16_9 ();
 sg13g2_decap_4 FILLER_16_18 ();
 sg13g2_fill_2 FILLER_16_35 ();
 sg13g2_fill_1 FILLER_16_37 ();
 sg13g2_decap_8 FILLER_16_62 ();
 sg13g2_fill_2 FILLER_16_69 ();
 sg13g2_decap_4 FILLER_16_90 ();
 sg13g2_fill_1 FILLER_16_110 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_4 FILLER_16_140 ();
 sg13g2_fill_1 FILLER_16_144 ();
 sg13g2_decap_4 FILLER_16_150 ();
 sg13g2_fill_2 FILLER_16_154 ();
 sg13g2_decap_4 FILLER_16_167 ();
 sg13g2_fill_1 FILLER_16_171 ();
 sg13g2_decap_4 FILLER_16_179 ();
 sg13g2_fill_1 FILLER_16_183 ();
 sg13g2_decap_8 FILLER_16_223 ();
 sg13g2_decap_4 FILLER_16_230 ();
 sg13g2_fill_2 FILLER_16_234 ();
 sg13g2_fill_2 FILLER_16_257 ();
 sg13g2_fill_1 FILLER_16_284 ();
 sg13g2_decap_4 FILLER_16_290 ();
 sg13g2_fill_1 FILLER_16_294 ();
 sg13g2_decap_4 FILLER_16_318 ();
 sg13g2_fill_1 FILLER_16_322 ();
 sg13g2_fill_1 FILLER_16_350 ();
 sg13g2_fill_1 FILLER_16_368 ();
 sg13g2_decap_4 FILLER_16_396 ();
 sg13g2_fill_1 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_41 ();
 sg13g2_fill_1 FILLER_17_48 ();
 sg13g2_fill_1 FILLER_17_69 ();
 sg13g2_fill_1 FILLER_17_79 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_decap_4 FILLER_17_95 ();
 sg13g2_fill_2 FILLER_17_99 ();
 sg13g2_decap_4 FILLER_17_114 ();
 sg13g2_fill_2 FILLER_17_118 ();
 sg13g2_fill_2 FILLER_17_138 ();
 sg13g2_fill_1 FILLER_17_140 ();
 sg13g2_decap_8 FILLER_17_154 ();
 sg13g2_fill_2 FILLER_17_161 ();
 sg13g2_fill_1 FILLER_17_169 ();
 sg13g2_fill_2 FILLER_17_176 ();
 sg13g2_fill_2 FILLER_17_197 ();
 sg13g2_fill_2 FILLER_17_206 ();
 sg13g2_fill_1 FILLER_17_208 ();
 sg13g2_fill_2 FILLER_17_214 ();
 sg13g2_fill_1 FILLER_17_216 ();
 sg13g2_decap_8 FILLER_17_223 ();
 sg13g2_fill_1 FILLER_17_230 ();
 sg13g2_fill_1 FILLER_17_244 ();
 sg13g2_decap_4 FILLER_17_254 ();
 sg13g2_fill_2 FILLER_17_258 ();
 sg13g2_decap_8 FILLER_17_272 ();
 sg13g2_fill_1 FILLER_17_279 ();
 sg13g2_fill_2 FILLER_17_295 ();
 sg13g2_decap_8 FILLER_17_309 ();
 sg13g2_fill_2 FILLER_17_316 ();
 sg13g2_fill_1 FILLER_17_318 ();
 sg13g2_decap_4 FILLER_17_337 ();
 sg13g2_decap_4 FILLER_17_347 ();
 sg13g2_fill_1 FILLER_17_364 ();
 sg13g2_fill_2 FILLER_17_378 ();
 sg13g2_fill_1 FILLER_17_380 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_2 FILLER_18_41 ();
 sg13g2_decap_4 FILLER_18_71 ();
 sg13g2_fill_2 FILLER_18_115 ();
 sg13g2_fill_1 FILLER_18_121 ();
 sg13g2_fill_2 FILLER_18_142 ();
 sg13g2_fill_1 FILLER_18_144 ();
 sg13g2_fill_2 FILLER_18_157 ();
 sg13g2_decap_4 FILLER_18_176 ();
 sg13g2_fill_2 FILLER_18_180 ();
 sg13g2_decap_4 FILLER_18_188 ();
 sg13g2_fill_2 FILLER_18_202 ();
 sg13g2_fill_1 FILLER_18_204 ();
 sg13g2_decap_4 FILLER_18_209 ();
 sg13g2_decap_4 FILLER_18_237 ();
 sg13g2_decap_4 FILLER_18_254 ();
 sg13g2_fill_1 FILLER_18_258 ();
 sg13g2_decap_8 FILLER_18_275 ();
 sg13g2_decap_4 FILLER_18_282 ();
 sg13g2_fill_1 FILLER_18_286 ();
 sg13g2_decap_4 FILLER_18_292 ();
 sg13g2_fill_1 FILLER_18_317 ();
 sg13g2_fill_2 FILLER_18_322 ();
 sg13g2_fill_1 FILLER_18_324 ();
 sg13g2_decap_4 FILLER_18_347 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_fill_1 FILLER_19_0 ();
 sg13g2_fill_2 FILLER_19_25 ();
 sg13g2_fill_1 FILLER_19_27 ();
 sg13g2_decap_4 FILLER_19_45 ();
 sg13g2_decap_4 FILLER_19_67 ();
 sg13g2_fill_1 FILLER_19_71 ();
 sg13g2_decap_8 FILLER_19_81 ();
 sg13g2_decap_8 FILLER_19_101 ();
 sg13g2_fill_1 FILLER_19_113 ();
 sg13g2_fill_1 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_4 FILLER_19_133 ();
 sg13g2_fill_1 FILLER_19_137 ();
 sg13g2_fill_2 FILLER_19_153 ();
 sg13g2_fill_1 FILLER_19_155 ();
 sg13g2_fill_2 FILLER_19_172 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_4 FILLER_19_203 ();
 sg13g2_fill_1 FILLER_19_207 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_fill_2 FILLER_19_231 ();
 sg13g2_decap_4 FILLER_19_238 ();
 sg13g2_fill_1 FILLER_19_247 ();
 sg13g2_decap_8 FILLER_19_257 ();
 sg13g2_fill_1 FILLER_19_276 ();
 sg13g2_decap_8 FILLER_19_313 ();
 sg13g2_fill_1 FILLER_19_320 ();
 sg13g2_decap_8 FILLER_19_347 ();
 sg13g2_decap_8 FILLER_19_372 ();
 sg13g2_decap_4 FILLER_19_379 ();
 sg13g2_fill_2 FILLER_20_0 ();
 sg13g2_fill_1 FILLER_20_2 ();
 sg13g2_fill_2 FILLER_20_7 ();
 sg13g2_fill_2 FILLER_20_35 ();
 sg13g2_decap_8 FILLER_20_41 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_fill_2 FILLER_20_55 ();
 sg13g2_decap_4 FILLER_20_63 ();
 sg13g2_fill_1 FILLER_20_67 ();
 sg13g2_fill_1 FILLER_20_73 ();
 sg13g2_fill_2 FILLER_20_85 ();
 sg13g2_fill_1 FILLER_20_87 ();
 sg13g2_fill_2 FILLER_20_97 ();
 sg13g2_fill_1 FILLER_20_99 ();
 sg13g2_fill_1 FILLER_20_111 ();
 sg13g2_fill_1 FILLER_20_129 ();
 sg13g2_fill_2 FILLER_20_180 ();
 sg13g2_fill_1 FILLER_20_182 ();
 sg13g2_decap_4 FILLER_20_189 ();
 sg13g2_fill_2 FILLER_20_221 ();
 sg13g2_decap_4 FILLER_20_227 ();
 sg13g2_decap_8 FILLER_20_254 ();
 sg13g2_fill_2 FILLER_20_261 ();
 sg13g2_fill_1 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_fill_2 FILLER_20_291 ();
 sg13g2_fill_1 FILLER_20_293 ();
 sg13g2_fill_2 FILLER_20_303 ();
 sg13g2_fill_1 FILLER_20_305 ();
 sg13g2_fill_2 FILLER_20_323 ();
 sg13g2_fill_1 FILLER_20_325 ();
 sg13g2_decap_8 FILLER_20_343 ();
 sg13g2_fill_2 FILLER_20_350 ();
 sg13g2_fill_1 FILLER_20_352 ();
 sg13g2_decap_4 FILLER_20_375 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_fill_2 FILLER_21_7 ();
 sg13g2_fill_1 FILLER_21_31 ();
 sg13g2_fill_2 FILLER_21_45 ();
 sg13g2_decap_8 FILLER_21_65 ();
 sg13g2_fill_2 FILLER_21_72 ();
 sg13g2_decap_4 FILLER_21_92 ();
 sg13g2_fill_1 FILLER_21_96 ();
 sg13g2_decap_8 FILLER_21_120 ();
 sg13g2_fill_1 FILLER_21_127 ();
 sg13g2_decap_8 FILLER_21_137 ();
 sg13g2_fill_2 FILLER_21_144 ();
 sg13g2_decap_8 FILLER_21_151 ();
 sg13g2_decap_4 FILLER_21_171 ();
 sg13g2_fill_2 FILLER_21_195 ();
 sg13g2_fill_1 FILLER_21_197 ();
 sg13g2_decap_4 FILLER_21_248 ();
 sg13g2_fill_1 FILLER_21_268 ();
 sg13g2_fill_1 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_289 ();
 sg13g2_decap_8 FILLER_21_313 ();
 sg13g2_decap_4 FILLER_21_320 ();
 sg13g2_fill_2 FILLER_21_324 ();
 sg13g2_decap_4 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_344 ();
 sg13g2_decap_4 FILLER_21_361 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_7 ();
 sg13g2_fill_2 FILLER_22_14 ();
 sg13g2_fill_1 FILLER_22_16 ();
 sg13g2_fill_1 FILLER_22_24 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_4 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_68 ();
 sg13g2_decap_4 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_97 ();
 sg13g2_decap_8 FILLER_22_121 ();
 sg13g2_fill_2 FILLER_22_140 ();
 sg13g2_fill_1 FILLER_22_142 ();
 sg13g2_fill_1 FILLER_22_161 ();
 sg13g2_fill_2 FILLER_22_167 ();
 sg13g2_fill_1 FILLER_22_169 ();
 sg13g2_decap_4 FILLER_22_180 ();
 sg13g2_fill_2 FILLER_22_184 ();
 sg13g2_fill_2 FILLER_22_199 ();
 sg13g2_fill_1 FILLER_22_201 ();
 sg13g2_decap_8 FILLER_22_218 ();
 sg13g2_decap_4 FILLER_22_233 ();
 sg13g2_decap_8 FILLER_22_241 ();
 sg13g2_decap_8 FILLER_22_248 ();
 sg13g2_fill_1 FILLER_22_255 ();
 sg13g2_decap_8 FILLER_22_274 ();
 sg13g2_decap_8 FILLER_22_287 ();
 sg13g2_fill_2 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_301 ();
 sg13g2_fill_1 FILLER_22_315 ();
 sg13g2_fill_1 FILLER_22_378 ();
 sg13g2_fill_2 FILLER_22_406 ();
 sg13g2_fill_1 FILLER_22_408 ();
 sg13g2_fill_2 FILLER_23_0 ();
 sg13g2_decap_4 FILLER_23_30 ();
 sg13g2_fill_2 FILLER_23_34 ();
 sg13g2_decap_4 FILLER_23_50 ();
 sg13g2_decap_4 FILLER_23_76 ();
 sg13g2_fill_1 FILLER_23_96 ();
 sg13g2_fill_2 FILLER_23_101 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_4 FILLER_23_126 ();
 sg13g2_decap_4 FILLER_23_138 ();
 sg13g2_fill_1 FILLER_23_142 ();
 sg13g2_fill_2 FILLER_23_148 ();
 sg13g2_fill_1 FILLER_23_150 ();
 sg13g2_decap_8 FILLER_23_156 ();
 sg13g2_decap_8 FILLER_23_163 ();
 sg13g2_decap_4 FILLER_23_170 ();
 sg13g2_fill_1 FILLER_23_174 ();
 sg13g2_fill_1 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_194 ();
 sg13g2_fill_2 FILLER_23_199 ();
 sg13g2_fill_2 FILLER_23_218 ();
 sg13g2_decap_4 FILLER_23_291 ();
 sg13g2_fill_1 FILLER_23_295 ();
 sg13g2_decap_4 FILLER_23_324 ();
 sg13g2_fill_2 FILLER_23_328 ();
 sg13g2_fill_1 FILLER_23_344 ();
 sg13g2_fill_2 FILLER_23_350 ();
 sg13g2_fill_1 FILLER_23_352 ();
 sg13g2_fill_2 FILLER_23_364 ();
 sg13g2_fill_1 FILLER_23_366 ();
 sg13g2_fill_1 FILLER_23_380 ();
 sg13g2_fill_2 FILLER_23_389 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_4 FILLER_24_11 ();
 sg13g2_fill_2 FILLER_24_15 ();
 sg13g2_fill_1 FILLER_24_22 ();
 sg13g2_fill_1 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_38 ();
 sg13g2_decap_4 FILLER_24_45 ();
 sg13g2_fill_1 FILLER_24_49 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_4 FILLER_24_79 ();
 sg13g2_fill_1 FILLER_24_83 ();
 sg13g2_fill_1 FILLER_24_102 ();
 sg13g2_decap_4 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_118 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_decap_4 FILLER_24_136 ();
 sg13g2_fill_1 FILLER_24_161 ();
 sg13g2_fill_1 FILLER_24_166 ();
 sg13g2_fill_1 FILLER_24_190 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_decap_4 FILLER_24_211 ();
 sg13g2_decap_8 FILLER_24_219 ();
 sg13g2_decap_8 FILLER_24_232 ();
 sg13g2_fill_2 FILLER_24_244 ();
 sg13g2_fill_2 FILLER_24_250 ();
 sg13g2_fill_1 FILLER_24_252 ();
 sg13g2_fill_1 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_261 ();
 sg13g2_decap_4 FILLER_24_284 ();
 sg13g2_fill_2 FILLER_24_288 ();
 sg13g2_decap_8 FILLER_24_294 ();
 sg13g2_fill_2 FILLER_24_301 ();
 sg13g2_fill_2 FILLER_24_315 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_340 ();
 sg13g2_fill_1 FILLER_24_346 ();
 sg13g2_fill_2 FILLER_24_373 ();
 sg13g2_fill_1 FILLER_24_380 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_13 ();
 sg13g2_decap_4 FILLER_25_20 ();
 sg13g2_fill_1 FILLER_25_24 ();
 sg13g2_decap_4 FILLER_25_48 ();
 sg13g2_fill_1 FILLER_25_52 ();
 sg13g2_fill_2 FILLER_25_63 ();
 sg13g2_fill_1 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_95 ();
 sg13g2_fill_2 FILLER_25_102 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_decap_8 FILLER_25_151 ();
 sg13g2_decap_8 FILLER_25_171 ();
 sg13g2_fill_2 FILLER_25_178 ();
 sg13g2_fill_1 FILLER_25_180 ();
 sg13g2_decap_8 FILLER_25_186 ();
 sg13g2_fill_1 FILLER_25_198 ();
 sg13g2_decap_8 FILLER_25_209 ();
 sg13g2_fill_1 FILLER_25_251 ();
 sg13g2_fill_2 FILLER_25_283 ();
 sg13g2_fill_2 FILLER_25_291 ();
 sg13g2_fill_1 FILLER_25_314 ();
 sg13g2_fill_2 FILLER_25_331 ();
 sg13g2_decap_4 FILLER_25_339 ();
 sg13g2_fill_1 FILLER_25_343 ();
 sg13g2_fill_1 FILLER_25_350 ();
 sg13g2_decap_4 FILLER_25_364 ();
 sg13g2_decap_4 FILLER_25_390 ();
 sg13g2_fill_2 FILLER_25_394 ();
 sg13g2_decap_8 FILLER_26_52 ();
 sg13g2_fill_1 FILLER_26_59 ();
 sg13g2_decap_8 FILLER_26_78 ();
 sg13g2_fill_2 FILLER_26_85 ();
 sg13g2_fill_1 FILLER_26_87 ();
 sg13g2_fill_2 FILLER_26_114 ();
 sg13g2_fill_1 FILLER_26_116 ();
 sg13g2_fill_1 FILLER_26_121 ();
 sg13g2_decap_4 FILLER_26_138 ();
 sg13g2_decap_4 FILLER_26_153 ();
 sg13g2_fill_1 FILLER_26_157 ();
 sg13g2_fill_1 FILLER_26_167 ();
 sg13g2_decap_8 FILLER_26_206 ();
 sg13g2_decap_8 FILLER_26_213 ();
 sg13g2_fill_2 FILLER_26_220 ();
 sg13g2_decap_8 FILLER_26_232 ();
 sg13g2_decap_4 FILLER_26_251 ();
 sg13g2_fill_2 FILLER_26_255 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_1 FILLER_26_263 ();
 sg13g2_decap_4 FILLER_26_268 ();
 sg13g2_decap_8 FILLER_26_276 ();
 sg13g2_decap_8 FILLER_26_283 ();
 sg13g2_fill_2 FILLER_26_309 ();
 sg13g2_fill_2 FILLER_26_316 ();
 sg13g2_fill_1 FILLER_26_345 ();
 sg13g2_decap_4 FILLER_26_363 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_fill_1 FILLER_26_379 ();
 sg13g2_fill_1 FILLER_26_408 ();
 sg13g2_decap_4 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_4 ();
 sg13g2_fill_2 FILLER_27_33 ();
 sg13g2_fill_1 FILLER_27_35 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_decap_8 FILLER_27_53 ();
 sg13g2_decap_4 FILLER_27_60 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_78 ();
 sg13g2_fill_1 FILLER_27_114 ();
 sg13g2_decap_8 FILLER_27_147 ();
 sg13g2_decap_4 FILLER_27_154 ();
 sg13g2_fill_2 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_173 ();
 sg13g2_decap_8 FILLER_27_180 ();
 sg13g2_fill_2 FILLER_27_187 ();
 sg13g2_fill_1 FILLER_27_189 ();
 sg13g2_fill_2 FILLER_27_205 ();
 sg13g2_decap_4 FILLER_27_213 ();
 sg13g2_fill_1 FILLER_27_237 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_decap_8 FILLER_27_273 ();
 sg13g2_decap_8 FILLER_27_287 ();
 sg13g2_decap_8 FILLER_27_299 ();
 sg13g2_fill_1 FILLER_27_345 ();
 sg13g2_fill_2 FILLER_27_351 ();
 sg13g2_fill_2 FILLER_27_358 ();
 sg13g2_fill_1 FILLER_27_360 ();
 sg13g2_fill_2 FILLER_27_371 ();
 sg13g2_fill_1 FILLER_27_373 ();
 sg13g2_decap_4 FILLER_27_379 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_7 ();
 sg13g2_fill_1 FILLER_28_9 ();
 sg13g2_decap_4 FILLER_28_14 ();
 sg13g2_fill_2 FILLER_28_18 ();
 sg13g2_fill_2 FILLER_28_65 ();
 sg13g2_fill_1 FILLER_28_67 ();
 sg13g2_fill_2 FILLER_28_77 ();
 sg13g2_fill_1 FILLER_28_79 ();
 sg13g2_fill_2 FILLER_28_97 ();
 sg13g2_fill_1 FILLER_28_99 ();
 sg13g2_decap_4 FILLER_28_105 ();
 sg13g2_fill_1 FILLER_28_109 ();
 sg13g2_decap_4 FILLER_28_119 ();
 sg13g2_fill_1 FILLER_28_123 ();
 sg13g2_fill_2 FILLER_28_134 ();
 sg13g2_fill_1 FILLER_28_136 ();
 sg13g2_fill_1 FILLER_28_162 ();
 sg13g2_fill_1 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_185 ();
 sg13g2_fill_1 FILLER_28_203 ();
 sg13g2_fill_2 FILLER_28_209 ();
 sg13g2_fill_1 FILLER_28_211 ();
 sg13g2_decap_8 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_247 ();
 sg13g2_fill_2 FILLER_28_269 ();
 sg13g2_fill_1 FILLER_28_271 ();
 sg13g2_fill_2 FILLER_28_304 ();
 sg13g2_fill_1 FILLER_28_312 ();
 sg13g2_fill_1 FILLER_28_324 ();
 sg13g2_fill_2 FILLER_28_366 ();
 sg13g2_fill_1 FILLER_28_368 ();
 sg13g2_fill_1 FILLER_28_373 ();
 sg13g2_fill_1 FILLER_28_392 ();
 sg13g2_fill_2 FILLER_28_406 ();
 sg13g2_fill_1 FILLER_28_408 ();
 sg13g2_fill_2 FILLER_29_32 ();
 sg13g2_fill_1 FILLER_29_34 ();
 sg13g2_fill_2 FILLER_29_44 ();
 sg13g2_fill_2 FILLER_29_59 ();
 sg13g2_fill_1 FILLER_29_61 ();
 sg13g2_decap_4 FILLER_29_68 ();
 sg13g2_decap_4 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_93 ();
 sg13g2_fill_1 FILLER_29_127 ();
 sg13g2_decap_8 FILLER_29_142 ();
 sg13g2_fill_2 FILLER_29_149 ();
 sg13g2_fill_1 FILLER_29_151 ();
 sg13g2_decap_4 FILLER_29_173 ();
 sg13g2_fill_2 FILLER_29_177 ();
 sg13g2_fill_2 FILLER_29_191 ();
 sg13g2_fill_2 FILLER_29_219 ();
 sg13g2_decap_4 FILLER_29_234 ();
 sg13g2_fill_1 FILLER_29_238 ();
 sg13g2_decap_8 FILLER_29_251 ();
 sg13g2_decap_4 FILLER_29_264 ();
 sg13g2_decap_4 FILLER_29_273 ();
 sg13g2_fill_2 FILLER_29_277 ();
 sg13g2_decap_4 FILLER_29_287 ();
 sg13g2_fill_2 FILLER_29_291 ();
 sg13g2_fill_1 FILLER_29_297 ();
 sg13g2_fill_1 FILLER_29_304 ();
 sg13g2_fill_2 FILLER_29_324 ();
 sg13g2_fill_1 FILLER_29_348 ();
 sg13g2_fill_1 FILLER_29_355 ();
 sg13g2_fill_2 FILLER_29_362 ();
 sg13g2_fill_1 FILLER_29_364 ();
 sg13g2_fill_2 FILLER_29_369 ();
 sg13g2_fill_1 FILLER_29_371 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_fill_1 FILLER_30_4 ();
 sg13g2_decap_4 FILLER_30_33 ();
 sg13g2_fill_2 FILLER_30_46 ();
 sg13g2_fill_1 FILLER_30_48 ();
 sg13g2_fill_1 FILLER_30_62 ();
 sg13g2_decap_4 FILLER_30_83 ();
 sg13g2_fill_2 FILLER_30_87 ();
 sg13g2_fill_2 FILLER_30_99 ();
 sg13g2_fill_1 FILLER_30_101 ();
 sg13g2_decap_8 FILLER_30_144 ();
 sg13g2_fill_1 FILLER_30_151 ();
 sg13g2_decap_4 FILLER_30_165 ();
 sg13g2_fill_2 FILLER_30_169 ();
 sg13g2_decap_4 FILLER_30_188 ();
 sg13g2_fill_1 FILLER_30_192 ();
 sg13g2_decap_8 FILLER_30_198 ();
 sg13g2_fill_2 FILLER_30_223 ();
 sg13g2_fill_2 FILLER_30_240 ();
 sg13g2_fill_2 FILLER_30_258 ();
 sg13g2_fill_1 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_288 ();
 sg13g2_fill_1 FILLER_30_306 ();
 sg13g2_fill_2 FILLER_30_318 ();
 sg13g2_decap_4 FILLER_30_328 ();
 sg13g2_fill_1 FILLER_30_332 ();
 sg13g2_decap_8 FILLER_30_341 ();
 sg13g2_fill_1 FILLER_30_348 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_368 ();
 sg13g2_fill_2 FILLER_30_397 ();
 sg13g2_fill_1 FILLER_30_408 ();
 sg13g2_decap_4 FILLER_31_0 ();
 sg13g2_fill_2 FILLER_31_4 ();
 sg13g2_fill_1 FILLER_31_14 ();
 sg13g2_fill_2 FILLER_31_32 ();
 sg13g2_fill_1 FILLER_31_34 ();
 sg13g2_decap_8 FILLER_31_78 ();
 sg13g2_decap_4 FILLER_31_85 ();
 sg13g2_fill_2 FILLER_31_107 ();
 sg13g2_decap_4 FILLER_31_139 ();
 sg13g2_fill_2 FILLER_31_143 ();
 sg13g2_fill_2 FILLER_31_156 ();
 sg13g2_decap_4 FILLER_31_164 ();
 sg13g2_fill_2 FILLER_31_176 ();
 sg13g2_fill_1 FILLER_31_195 ();
 sg13g2_fill_1 FILLER_31_215 ();
 sg13g2_fill_2 FILLER_31_226 ();
 sg13g2_decap_8 FILLER_31_233 ();
 sg13g2_fill_2 FILLER_31_240 ();
 sg13g2_decap_8 FILLER_31_265 ();
 sg13g2_fill_2 FILLER_31_287 ();
 sg13g2_fill_1 FILLER_31_289 ();
 sg13g2_decap_8 FILLER_31_300 ();
 sg13g2_decap_8 FILLER_31_307 ();
 sg13g2_fill_1 FILLER_31_314 ();
 sg13g2_decap_4 FILLER_31_323 ();
 sg13g2_fill_2 FILLER_31_336 ();
 sg13g2_fill_1 FILLER_31_351 ();
 sg13g2_fill_1 FILLER_31_362 ();
 sg13g2_fill_2 FILLER_32_0 ();
 sg13g2_fill_2 FILLER_32_15 ();
 sg13g2_decap_4 FILLER_32_29 ();
 sg13g2_fill_1 FILLER_32_33 ();
 sg13g2_decap_4 FILLER_32_47 ();
 sg13g2_decap_4 FILLER_32_58 ();
 sg13g2_fill_2 FILLER_32_74 ();
 sg13g2_fill_1 FILLER_32_76 ();
 sg13g2_decap_4 FILLER_32_89 ();
 sg13g2_fill_1 FILLER_32_98 ();
 sg13g2_fill_2 FILLER_32_109 ();
 sg13g2_fill_1 FILLER_32_111 ();
 sg13g2_decap_4 FILLER_32_116 ();
 sg13g2_fill_1 FILLER_32_120 ();
 sg13g2_fill_1 FILLER_32_168 ();
 sg13g2_fill_2 FILLER_32_179 ();
 sg13g2_fill_1 FILLER_32_181 ();
 sg13g2_fill_2 FILLER_32_190 ();
 sg13g2_fill_1 FILLER_32_192 ();
 sg13g2_decap_4 FILLER_32_209 ();
 sg13g2_fill_2 FILLER_32_213 ();
 sg13g2_decap_8 FILLER_32_224 ();
 sg13g2_decap_4 FILLER_32_231 ();
 sg13g2_fill_1 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_fill_2 FILLER_32_270 ();
 sg13g2_fill_1 FILLER_32_272 ();
 sg13g2_decap_4 FILLER_32_282 ();
 sg13g2_fill_2 FILLER_32_309 ();
 sg13g2_decap_4 FILLER_32_345 ();
 sg13g2_fill_2 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_366 ();
 sg13g2_fill_1 FILLER_32_394 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_11 ();
 sg13g2_fill_2 FILLER_33_18 ();
 sg13g2_decap_4 FILLER_33_48 ();
 sg13g2_fill_2 FILLER_33_64 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_fill_1 FILLER_33_93 ();
 sg13g2_decap_8 FILLER_33_99 ();
 sg13g2_decap_8 FILLER_33_106 ();
 sg13g2_fill_1 FILLER_33_113 ();
 sg13g2_decap_4 FILLER_33_123 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_150 ();
 sg13g2_fill_2 FILLER_33_169 ();
 sg13g2_fill_2 FILLER_33_176 ();
 sg13g2_fill_2 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_238 ();
 sg13g2_fill_2 FILLER_33_248 ();
 sg13g2_fill_1 FILLER_33_250 ();
 sg13g2_decap_4 FILLER_33_262 ();
 sg13g2_fill_2 FILLER_33_281 ();
 sg13g2_fill_1 FILLER_33_283 ();
 sg13g2_fill_2 FILLER_33_293 ();
 sg13g2_fill_1 FILLER_33_295 ();
 sg13g2_decap_4 FILLER_33_310 ();
 sg13g2_fill_2 FILLER_33_314 ();
 sg13g2_decap_4 FILLER_33_323 ();
 sg13g2_fill_2 FILLER_33_327 ();
 sg13g2_decap_8 FILLER_33_338 ();
 sg13g2_decap_4 FILLER_33_345 ();
 sg13g2_fill_1 FILLER_33_354 ();
 sg13g2_decap_4 FILLER_33_361 ();
 sg13g2_fill_2 FILLER_33_365 ();
 sg13g2_decap_8 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_7 ();
 sg13g2_decap_8 FILLER_34_12 ();
 sg13g2_decap_4 FILLER_34_19 ();
 sg13g2_fill_2 FILLER_34_23 ();
 sg13g2_fill_2 FILLER_34_43 ();
 sg13g2_decap_4 FILLER_34_59 ();
 sg13g2_decap_8 FILLER_34_68 ();
 sg13g2_decap_8 FILLER_34_75 ();
 sg13g2_fill_1 FILLER_34_82 ();
 sg13g2_fill_2 FILLER_34_102 ();
 sg13g2_fill_1 FILLER_34_104 ();
 sg13g2_decap_8 FILLER_34_122 ();
 sg13g2_decap_8 FILLER_34_129 ();
 sg13g2_decap_4 FILLER_34_136 ();
 sg13g2_fill_2 FILLER_34_140 ();
 sg13g2_fill_1 FILLER_34_157 ();
 sg13g2_fill_1 FILLER_34_176 ();
 sg13g2_fill_2 FILLER_34_219 ();
 sg13g2_decap_4 FILLER_34_256 ();
 sg13g2_fill_1 FILLER_34_260 ();
 sg13g2_fill_2 FILLER_34_292 ();
 sg13g2_fill_2 FILLER_34_308 ();
 sg13g2_decap_4 FILLER_34_324 ();
 sg13g2_fill_1 FILLER_34_343 ();
 sg13g2_fill_2 FILLER_34_362 ();
 sg13g2_fill_1 FILLER_34_378 ();
 sg13g2_fill_2 FILLER_34_389 ();
 sg13g2_fill_1 FILLER_34_391 ();
 sg13g2_fill_2 FILLER_35_0 ();
 sg13g2_fill_1 FILLER_35_2 ();
 sg13g2_decap_4 FILLER_35_92 ();
 sg13g2_decap_4 FILLER_35_110 ();
 sg13g2_decap_4 FILLER_35_134 ();
 sg13g2_fill_1 FILLER_35_167 ();
 sg13g2_fill_2 FILLER_35_177 ();
 sg13g2_fill_2 FILLER_35_218 ();
 sg13g2_fill_1 FILLER_35_220 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_256 ();
 sg13g2_fill_2 FILLER_35_266 ();
 sg13g2_decap_4 FILLER_35_282 ();
 sg13g2_fill_2 FILLER_35_294 ();
 sg13g2_fill_2 FILLER_35_303 ();
 sg13g2_fill_1 FILLER_35_305 ();
 sg13g2_fill_1 FILLER_35_313 ();
 sg13g2_decap_4 FILLER_35_326 ();
 sg13g2_fill_1 FILLER_35_330 ();
 sg13g2_fill_2 FILLER_35_345 ();
 sg13g2_fill_2 FILLER_35_379 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_39 ();
 sg13g2_decap_4 FILLER_36_50 ();
 sg13g2_decap_4 FILLER_36_72 ();
 sg13g2_fill_1 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_95 ();
 sg13g2_decap_4 FILLER_36_127 ();
 sg13g2_fill_1 FILLER_36_169 ();
 sg13g2_decap_4 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_190 ();
 sg13g2_decap_8 FILLER_36_205 ();
 sg13g2_decap_8 FILLER_36_212 ();
 sg13g2_decap_8 FILLER_36_219 ();
 sg13g2_fill_2 FILLER_36_226 ();
 sg13g2_fill_1 FILLER_36_228 ();
 sg13g2_fill_2 FILLER_36_274 ();
 sg13g2_fill_1 FILLER_36_276 ();
 sg13g2_fill_2 FILLER_36_288 ();
 sg13g2_fill_1 FILLER_36_312 ();
 sg13g2_fill_2 FILLER_36_339 ();
 sg13g2_fill_1 FILLER_36_391 ();
 sg13g2_fill_2 FILLER_36_406 ();
 sg13g2_fill_1 FILLER_36_408 ();
 sg13g2_fill_1 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_74 ();
 sg13g2_fill_1 FILLER_37_80 ();
 sg13g2_fill_2 FILLER_37_96 ();
 sg13g2_fill_1 FILLER_37_98 ();
 sg13g2_decap_8 FILLER_37_135 ();
 sg13g2_decap_4 FILLER_37_142 ();
 sg13g2_fill_1 FILLER_37_146 ();
 sg13g2_decap_4 FILLER_37_167 ();
 sg13g2_fill_2 FILLER_37_171 ();
 sg13g2_decap_8 FILLER_37_177 ();
 sg13g2_decap_8 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_191 ();
 sg13g2_decap_4 FILLER_37_223 ();
 sg13g2_fill_1 FILLER_37_227 ();
 sg13g2_fill_1 FILLER_37_254 ();
 sg13g2_fill_1 FILLER_37_293 ();
 sg13g2_fill_1 FILLER_37_303 ();
 sg13g2_fill_1 FILLER_37_335 ();
 sg13g2_fill_2 FILLER_37_349 ();
 sg13g2_fill_1 FILLER_37_351 ();
 sg13g2_fill_2 FILLER_37_378 ();
 sg13g2_fill_1 FILLER_37_380 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_2 FILLER_38_47 ();
 sg13g2_fill_2 FILLER_38_58 ();
 sg13g2_fill_2 FILLER_38_109 ();
 sg13g2_fill_1 FILLER_38_111 ();
 sg13g2_decap_8 FILLER_38_148 ();
 sg13g2_decap_8 FILLER_38_155 ();
 sg13g2_decap_4 FILLER_38_162 ();
 sg13g2_fill_2 FILLER_38_166 ();
 sg13g2_fill_1 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_201 ();
 sg13g2_fill_1 FILLER_38_319 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
endmodule
