module tt_um_rebeccargb_intercal_alu (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire clknet_0_clk;
 wire \a[0] ;
 wire \a[10] ;
 wire \a[11] ;
 wire \a[12] ;
 wire \a[13] ;
 wire \a[14] ;
 wire \a[15] ;
 wire \a[16] ;
 wire \a[17] ;
 wire \a[18] ;
 wire \a[19] ;
 wire \a[1] ;
 wire \a[20] ;
 wire \a[21] ;
 wire \a[22] ;
 wire \a[23] ;
 wire \a[24] ;
 wire \a[25] ;
 wire \a[26] ;
 wire \a[27] ;
 wire \a[28] ;
 wire \a[29] ;
 wire \a[2] ;
 wire \a[30] ;
 wire \a[31] ;
 wire \a[3] ;
 wire \a[4] ;
 wire \a[5] ;
 wire \a[6] ;
 wire \a[7] ;
 wire \a[8] ;
 wire \a[9] ;
 wire \ayayayayayaya.b[0] ;
 wire \ayayayayayaya.b[10] ;
 wire \ayayayayayaya.b[11] ;
 wire \ayayayayayaya.b[12] ;
 wire \ayayayayayaya.b[13] ;
 wire \ayayayayayaya.b[14] ;
 wire \ayayayayayaya.b[15] ;
 wire \ayayayayayaya.b[16] ;
 wire \ayayayayayaya.b[17] ;
 wire \ayayayayayaya.b[18] ;
 wire \ayayayayayaya.b[19] ;
 wire \ayayayayayaya.b[1] ;
 wire \ayayayayayaya.b[20] ;
 wire \ayayayayayaya.b[21] ;
 wire \ayayayayayaya.b[22] ;
 wire \ayayayayayaya.b[23] ;
 wire \ayayayayayaya.b[24] ;
 wire \ayayayayayaya.b[25] ;
 wire \ayayayayayaya.b[26] ;
 wire \ayayayayayaya.b[27] ;
 wire \ayayayayayaya.b[28] ;
 wire \ayayayayayaya.b[29] ;
 wire \ayayayayayaya.b[2] ;
 wire \ayayayayayaya.b[30] ;
 wire \ayayayayayaya.b[31] ;
 wire \ayayayayayaya.b[3] ;
 wire \ayayayayayaya.b[4] ;
 wire \ayayayayayaya.b[5] ;
 wire \ayayayayayaya.b[6] ;
 wire \ayayayayayaya.b[7] ;
 wire \ayayayayayaya.b[8] ;
 wire \ayayayayayaya.b[9] ;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;

 sg13g2_inv_4 _1742_ (.A(net843),
    .Y(_0600_));
 sg13g2_inv_4 _1743_ (.A(net847),
    .Y(_0611_));
 sg13g2_inv_2 _1744_ (.Y(_0621_),
    .A(net81));
 sg13g2_inv_1 _1745_ (.Y(_0632_),
    .A(net100));
 sg13g2_inv_2 _1746_ (.Y(_0643_),
    .A(net82));
 sg13g2_inv_2 _1747_ (.Y(_0654_),
    .A(net101));
 sg13g2_inv_1 _1748_ (.Y(_0665_),
    .A(net829));
 sg13g2_inv_1 _1749_ (.Y(_0676_),
    .A(net91));
 sg13g2_inv_2 _1750_ (.Y(_0686_),
    .A(net87));
 sg13g2_inv_2 _1751_ (.Y(_0697_),
    .A(net111));
 sg13g2_inv_2 _1752_ (.Y(_0708_),
    .A(net716));
 sg13g2_inv_1 _1753_ (.Y(_0719_),
    .A(net717));
 sg13g2_inv_1 _1754_ (.Y(_0730_),
    .A(net718));
 sg13g2_inv_1 _1755_ (.Y(_0740_),
    .A(net719));
 sg13g2_inv_1 _1756_ (.Y(_0751_),
    .A(net721));
 sg13g2_inv_2 _1757_ (.Y(_0762_),
    .A(net723));
 sg13g2_inv_1 _1758_ (.Y(_0773_),
    .A(net726));
 sg13g2_inv_1 _1759_ (.Y(_0784_),
    .A(net727));
 sg13g2_inv_1 _1760_ (.Y(_0795_),
    .A(net729));
 sg13g2_inv_1 _1761_ (.Y(_0806_),
    .A(net732));
 sg13g2_inv_1 _1762_ (.Y(_0810_),
    .A(net735));
 sg13g2_inv_1 _1763_ (.Y(_0813_),
    .A(net739));
 sg13g2_inv_1 _1764_ (.Y(_0818_),
    .A(net743));
 sg13g2_inv_1 _1765_ (.Y(_0823_),
    .A(net747));
 sg13g2_inv_1 _1766_ (.Y(_0826_),
    .A(net750));
 sg13g2_inv_1 _1767_ (.Y(_0832_),
    .A(net755));
 sg13g2_inv_2 _1768_ (.Y(_0839_),
    .A(net760));
 sg13g2_inv_1 _1769_ (.Y(_0845_),
    .A(net765));
 sg13g2_inv_1 _1770_ (.Y(_0851_),
    .A(net770));
 sg13g2_inv_1 _1771_ (.Y(_0858_),
    .A(net774));
 sg13g2_inv_2 _1772_ (.Y(_0863_),
    .A(net780));
 sg13g2_inv_1 _1773_ (.Y(_0864_),
    .A(net786));
 sg13g2_inv_1 _1774_ (.Y(_0865_),
    .A(net793));
 sg13g2_inv_2 _1775_ (.Y(_0866_),
    .A(net800));
 sg13g2_inv_1 _1776_ (.Y(_0867_),
    .A(net807));
 sg13g2_inv_4 _1777_ (.A(net814),
    .Y(_0868_));
 sg13g2_inv_2 _1778_ (.Y(uio_oe[7]),
    .A(net4));
 sg13g2_nor2b_2 _1779_ (.A(net2),
    .B_N(net3),
    .Y(_0869_));
 sg13g2_and3_2 _1780_ (.X(_0870_),
    .A(net840),
    .B(net1),
    .C(_0869_));
 sg13g2_nand3_1 _1781_ (.B(net1),
    .C(_0869_),
    .A(net840),
    .Y(_0871_));
 sg13g2_and2_1 _1782_ (.A(net822),
    .B(_0870_),
    .X(_0872_));
 sg13g2_nand2_1 _1783_ (.Y(_0873_),
    .A(net822),
    .B(_0870_));
 sg13g2_and4_1 _1784_ (.A(\a[31] ),
    .B(\ayayayayayaya.b[31] ),
    .C(\ayayayayayaya.b[30] ),
    .D(\ayayayayayaya.b[29] ),
    .X(_0874_));
 sg13g2_a21oi_1 _1785_ (.A1(\a[31] ),
    .A2(\ayayayayayaya.b[31] ),
    .Y(_0875_),
    .B1(\ayayayayayaya.b[30] ));
 sg13g2_nor2b_1 _1786_ (.A(\a[30] ),
    .B_N(\ayayayayayaya.b[30] ),
    .Y(_0876_));
 sg13g2_and4_1 _1787_ (.A(net829),
    .B(\ayayayayayaya.b[31] ),
    .C(\ayayayayayaya.b[30] ),
    .D(_0676_),
    .X(_0877_));
 sg13g2_nor3_1 _1788_ (.A(_0676_),
    .B(_0875_),
    .C(_0876_),
    .Y(_0878_));
 sg13g2_nor3_1 _1789_ (.A(_0686_),
    .B(_0877_),
    .C(_0878_),
    .Y(_0879_));
 sg13g2_nor2_1 _1790_ (.A(\ayayayayayaya.b[28] ),
    .B(_0874_),
    .Y(_0880_));
 sg13g2_and2_1 _1791_ (.A(\ayayayayayaya.b[28] ),
    .B(_0874_),
    .X(_0881_));
 sg13g2_and2_1 _1792_ (.A(_0697_),
    .B(_0881_),
    .X(_0882_));
 sg13g2_nor3_1 _1793_ (.A(_0697_),
    .B(_0879_),
    .C(_0880_),
    .Y(_0883_));
 sg13g2_and2_1 _1794_ (.A(\a[29] ),
    .B(\ayayayayayaya.b[29] ),
    .X(_0884_));
 sg13g2_nor3_1 _1795_ (.A(\ayayayayayaya.b[29] ),
    .B(_0875_),
    .C(_0876_),
    .Y(_0885_));
 sg13g2_nor3_1 _1796_ (.A(_0686_),
    .B(_0884_),
    .C(_0885_),
    .Y(_0886_));
 sg13g2_nor3_1 _1797_ (.A(\ayayayayayaya.b[28] ),
    .B(_0877_),
    .C(_0878_),
    .Y(_0887_));
 sg13g2_nor3_1 _1798_ (.A(\ayayayayayaya.b[27] ),
    .B(_0879_),
    .C(_0880_),
    .Y(_0888_));
 sg13g2_nor3_1 _1799_ (.A(_0697_),
    .B(_0886_),
    .C(_0887_),
    .Y(_0889_));
 sg13g2_nor3_1 _1800_ (.A(_0708_),
    .B(_0888_),
    .C(_0889_),
    .Y(_0890_));
 sg13g2_nor3_1 _1801_ (.A(net716),
    .B(_0882_),
    .C(_0883_),
    .Y(_0891_));
 sg13g2_nor3_1 _1802_ (.A(_0708_),
    .B(_0882_),
    .C(_0883_),
    .Y(_0892_));
 sg13g2_a21oi_1 _1803_ (.A1(\ayayayayayaya.b[27] ),
    .A2(_0881_),
    .Y(_0893_),
    .B1(net716));
 sg13g2_nor3_1 _1804_ (.A(net717),
    .B(_0892_),
    .C(_0893_),
    .Y(_0894_));
 sg13g2_nor3_1 _1805_ (.A(net715),
    .B(_0890_),
    .C(_0891_),
    .Y(_0895_));
 sg13g2_nor3_1 _1806_ (.A(\ayayayayayaya.b[28] ),
    .B(_0884_),
    .C(_0885_),
    .Y(_0896_));
 sg13g2_nor2_1 _1807_ (.A(\a[28] ),
    .B(_0686_),
    .Y(_0897_));
 sg13g2_nor3_1 _1808_ (.A(\ayayayayayaya.b[27] ),
    .B(_0886_),
    .C(_0887_),
    .Y(_0898_));
 sg13g2_nor3_1 _1809_ (.A(_0697_),
    .B(_0896_),
    .C(_0897_),
    .Y(_0899_));
 sg13g2_nor3_1 _1810_ (.A(_0708_),
    .B(_0898_),
    .C(_0899_),
    .Y(_0900_));
 sg13g2_nor3_1 _1811_ (.A(net716),
    .B(_0888_),
    .C(_0889_),
    .Y(_0901_));
 sg13g2_nor3_1 _1812_ (.A(net717),
    .B(_0890_),
    .C(_0891_),
    .Y(_0902_));
 sg13g2_nor3_1 _1813_ (.A(net715),
    .B(_0900_),
    .C(_0901_),
    .Y(_0903_));
 sg13g2_nor3_1 _1814_ (.A(net714),
    .B(_0902_),
    .C(_0903_),
    .Y(_0904_));
 sg13g2_nor3_1 _1815_ (.A(net718),
    .B(_0894_),
    .C(_0895_),
    .Y(_0905_));
 sg13g2_o21ai_1 _1816_ (.B1(_0697_),
    .Y(_0906_),
    .A1(_0896_),
    .A2(_0897_));
 sg13g2_nand2b_1 _1817_ (.Y(_0907_),
    .B(\ayayayayayaya.b[27] ),
    .A_N(\a[27] ));
 sg13g2_o21ai_1 _1818_ (.B1(_0708_),
    .Y(_0908_),
    .A1(_0898_),
    .A2(_0899_));
 sg13g2_nand3_1 _1819_ (.B(_0906_),
    .C(_0907_),
    .A(net716),
    .Y(_0909_));
 sg13g2_nand3_1 _1820_ (.B(_0908_),
    .C(_0909_),
    .A(net717),
    .Y(_0910_));
 sg13g2_o21ai_1 _1821_ (.B1(net715),
    .Y(_0911_),
    .A1(_0900_),
    .A2(_0901_));
 sg13g2_o21ai_1 _1822_ (.B1(net714),
    .Y(_0912_),
    .A1(_0902_),
    .A2(_0903_));
 sg13g2_nand3_1 _1823_ (.B(_0910_),
    .C(_0911_),
    .A(net718),
    .Y(_0913_));
 sg13g2_nand3_1 _1824_ (.B(_0912_),
    .C(_0913_),
    .A(net719),
    .Y(_0914_));
 sg13g2_o21ai_1 _1825_ (.B1(net713),
    .Y(_0915_),
    .A1(_0904_),
    .A2(_0905_));
 sg13g2_nand3_1 _1826_ (.B(net716),
    .C(_0881_),
    .A(\ayayayayayaya.b[27] ),
    .Y(_0916_));
 sg13g2_nor2_1 _1827_ (.A(\ayayayayayaya.b[25] ),
    .B(_0916_),
    .Y(_0917_));
 sg13g2_nor3_1 _1828_ (.A(net715),
    .B(_0892_),
    .C(_0893_),
    .Y(_0918_));
 sg13g2_nor3_1 _1829_ (.A(net714),
    .B(_0894_),
    .C(_0895_),
    .Y(_0919_));
 sg13g2_nor3_1 _1830_ (.A(\ayayayayayaya.b[24] ),
    .B(_0917_),
    .C(_0918_),
    .Y(_0920_));
 sg13g2_nor3_1 _1831_ (.A(net719),
    .B(_0919_),
    .C(_0920_),
    .Y(_0921_));
 sg13g2_nor3_1 _1832_ (.A(net713),
    .B(_0904_),
    .C(_0905_),
    .Y(_0922_));
 sg13g2_o21ai_1 _1833_ (.B1(net711),
    .Y(_0923_),
    .A1(_0921_),
    .A2(_0922_));
 sg13g2_nand3_1 _1834_ (.B(_0914_),
    .C(_0915_),
    .A(net721),
    .Y(_0924_));
 sg13g2_a21oi_1 _1835_ (.A1(_0906_),
    .A2(_0907_),
    .Y(_0925_),
    .B1(\ayayayayayaya.b[26] ));
 sg13g2_nor2_1 _1836_ (.A(\a[26] ),
    .B(_0708_),
    .Y(_0926_));
 sg13g2_o21ai_1 _1837_ (.B1(net717),
    .Y(_0927_),
    .A1(_0925_),
    .A2(_0926_));
 sg13g2_nand3_1 _1838_ (.B(_0908_),
    .C(_0909_),
    .A(net715),
    .Y(_0928_));
 sg13g2_nand3_1 _1839_ (.B(_0910_),
    .C(_0911_),
    .A(net714),
    .Y(_0929_));
 sg13g2_nand3_1 _1840_ (.B(_0927_),
    .C(_0928_),
    .A(net718),
    .Y(_0930_));
 sg13g2_nand3_1 _1841_ (.B(_0929_),
    .C(_0930_),
    .A(net719),
    .Y(_0931_));
 sg13g2_nand3_1 _1842_ (.B(_0912_),
    .C(_0913_),
    .A(net713),
    .Y(_0932_));
 sg13g2_nand3_1 _1843_ (.B(_0914_),
    .C(_0915_),
    .A(net711),
    .Y(_0933_));
 sg13g2_nand3_1 _1844_ (.B(_0931_),
    .C(_0932_),
    .A(net721),
    .Y(_0934_));
 sg13g2_nand3_1 _1845_ (.B(_0933_),
    .C(_0934_),
    .A(net723),
    .Y(_0935_));
 sg13g2_nand3_1 _1846_ (.B(_0923_),
    .C(_0924_),
    .A(net710),
    .Y(_0936_));
 sg13g2_nor2_1 _1847_ (.A(net715),
    .B(_0916_),
    .Y(_0937_));
 sg13g2_nor3_1 _1848_ (.A(net714),
    .B(_0917_),
    .C(_0918_),
    .Y(_0938_));
 sg13g2_nor2_1 _1849_ (.A(\ayayayayayaya.b[24] ),
    .B(_0937_),
    .Y(_0939_));
 sg13g2_nor3_1 _1850_ (.A(net719),
    .B(_0938_),
    .C(_0939_),
    .Y(_0940_));
 sg13g2_nor3_1 _1851_ (.A(net713),
    .B(_0919_),
    .C(_0920_),
    .Y(_0941_));
 sg13g2_nor3_1 _1852_ (.A(net711),
    .B(_0921_),
    .C(_0922_),
    .Y(_0942_));
 sg13g2_nor3_1 _1853_ (.A(net721),
    .B(_0940_),
    .C(_0941_),
    .Y(_0943_));
 sg13g2_nand3_1 _1854_ (.B(_0923_),
    .C(_0924_),
    .A(net723),
    .Y(_0944_));
 sg13g2_o21ai_1 _1855_ (.B1(net710),
    .Y(_0945_),
    .A1(_0942_),
    .A2(_0943_));
 sg13g2_nand3_1 _1856_ (.B(_0944_),
    .C(_0945_),
    .A(net709),
    .Y(_0946_));
 sg13g2_nand3_1 _1857_ (.B(_0935_),
    .C(_0936_),
    .A(net725),
    .Y(_0947_));
 sg13g2_o21ai_1 _1858_ (.B1(net715),
    .Y(_0948_),
    .A1(_0925_),
    .A2(_0926_));
 sg13g2_nand2b_1 _1859_ (.Y(_0949_),
    .B(net717),
    .A_N(\a[25] ));
 sg13g2_nand3_1 _1860_ (.B(_0927_),
    .C(_0928_),
    .A(net714),
    .Y(_0950_));
 sg13g2_nand3_1 _1861_ (.B(_0948_),
    .C(_0949_),
    .A(net718),
    .Y(_0951_));
 sg13g2_nand3_1 _1862_ (.B(_0950_),
    .C(_0951_),
    .A(net719),
    .Y(_0952_));
 sg13g2_nand3_1 _1863_ (.B(_0929_),
    .C(_0930_),
    .A(net713),
    .Y(_0953_));
 sg13g2_nand3_1 _1864_ (.B(_0931_),
    .C(_0932_),
    .A(net711),
    .Y(_0954_));
 sg13g2_nand3_1 _1865_ (.B(_0952_),
    .C(_0953_),
    .A(net721),
    .Y(_0955_));
 sg13g2_nand3_1 _1866_ (.B(_0954_),
    .C(_0955_),
    .A(net722),
    .Y(_0956_));
 sg13g2_nand3_1 _1867_ (.B(_0933_),
    .C(_0934_),
    .A(net710),
    .Y(_0957_));
 sg13g2_nand3_1 _1868_ (.B(_0935_),
    .C(_0936_),
    .A(net709),
    .Y(_0958_));
 sg13g2_nand3_1 _1869_ (.B(_0956_),
    .C(_0957_),
    .A(net725),
    .Y(_0959_));
 sg13g2_nand3_1 _1870_ (.B(_0958_),
    .C(_0959_),
    .A(net727),
    .Y(_0960_));
 sg13g2_nand3_1 _1871_ (.B(_0946_),
    .C(_0947_),
    .A(net706),
    .Y(_0961_));
 sg13g2_nor4_1 _1872_ (.A(_0719_),
    .B(_0730_),
    .C(net719),
    .D(_0916_),
    .Y(_0962_));
 sg13g2_nor3_1 _1873_ (.A(net713),
    .B(_0938_),
    .C(_0939_),
    .Y(_0963_));
 sg13g2_nor3_1 _1874_ (.A(net712),
    .B(_0940_),
    .C(_0941_),
    .Y(_0964_));
 sg13g2_nor3_1 _1875_ (.A(\ayayayayayaya.b[22] ),
    .B(_0962_),
    .C(_0963_),
    .Y(_0965_));
 sg13g2_nor3_1 _1876_ (.A(net722),
    .B(_0964_),
    .C(_0965_),
    .Y(_0966_));
 sg13g2_nor3_1 _1877_ (.A(_0762_),
    .B(_0942_),
    .C(_0943_),
    .Y(_0967_));
 sg13g2_o21ai_1 _1878_ (.B1(net709),
    .Y(_0968_),
    .A1(_0966_),
    .A2(_0967_));
 sg13g2_nand3_1 _1879_ (.B(_0944_),
    .C(_0945_),
    .A(net725),
    .Y(_0969_));
 sg13g2_nand3_1 _1880_ (.B(_0946_),
    .C(_0947_),
    .A(net727),
    .Y(_0970_));
 sg13g2_nand3_1 _1881_ (.B(_0968_),
    .C(_0969_),
    .A(net706),
    .Y(_0971_));
 sg13g2_nand3_1 _1882_ (.B(_0970_),
    .C(_0971_),
    .A(net704),
    .Y(_0972_));
 sg13g2_nand3_1 _1883_ (.B(_0960_),
    .C(_0961_),
    .A(net729),
    .Y(_0973_));
 sg13g2_a21oi_1 _1884_ (.A1(_0948_),
    .A2(_0949_),
    .Y(_0974_),
    .B1(net718));
 sg13g2_nor2_1 _1885_ (.A(\a[24] ),
    .B(net714),
    .Y(_0975_));
 sg13g2_o21ai_1 _1886_ (.B1(net719),
    .Y(_0976_),
    .A1(_0974_),
    .A2(_0975_));
 sg13g2_nand3_1 _1887_ (.B(_0950_),
    .C(_0951_),
    .A(net713),
    .Y(_0977_));
 sg13g2_nand3_1 _1888_ (.B(_0952_),
    .C(_0953_),
    .A(net711),
    .Y(_0978_));
 sg13g2_nand3_1 _1889_ (.B(_0976_),
    .C(_0977_),
    .A(\ayayayayayaya.b[22] ),
    .Y(_0979_));
 sg13g2_nand3_1 _1890_ (.B(_0978_),
    .C(_0979_),
    .A(net722),
    .Y(_0980_));
 sg13g2_nand3_1 _1891_ (.B(_0954_),
    .C(_0955_),
    .A(net710),
    .Y(_0981_));
 sg13g2_nand3_1 _1892_ (.B(_0956_),
    .C(_0957_),
    .A(net708),
    .Y(_0982_));
 sg13g2_nand3_1 _1893_ (.B(_0980_),
    .C(_0981_),
    .A(net725),
    .Y(_0983_));
 sg13g2_nand3_1 _1894_ (.B(_0982_),
    .C(_0983_),
    .A(net727),
    .Y(_0984_));
 sg13g2_nand3_1 _1895_ (.B(_0958_),
    .C(_0959_),
    .A(net706),
    .Y(_0985_));
 sg13g2_nand3_1 _1896_ (.B(_0960_),
    .C(_0961_),
    .A(net704),
    .Y(_0986_));
 sg13g2_nand3_1 _1897_ (.B(_0984_),
    .C(_0985_),
    .A(net729),
    .Y(_0987_));
 sg13g2_nand3_1 _1898_ (.B(_0986_),
    .C(_0987_),
    .A(net732),
    .Y(_0988_));
 sg13g2_nand3_1 _1899_ (.B(_0972_),
    .C(_0973_),
    .A(net702),
    .Y(_0989_));
 sg13g2_nand3_1 _1900_ (.B(net720),
    .C(_0937_),
    .A(\ayayayayayaya.b[24] ),
    .Y(_0990_));
 sg13g2_nor3_1 _1901_ (.A(net712),
    .B(_0962_),
    .C(_0963_),
    .Y(_0991_));
 sg13g2_and2_1 _1902_ (.A(net712),
    .B(_0990_),
    .X(_0992_));
 sg13g2_nor3_1 _1903_ (.A(net723),
    .B(_0991_),
    .C(_0992_),
    .Y(_0993_));
 sg13g2_nor3_1 _1904_ (.A(_0762_),
    .B(_0964_),
    .C(_0965_),
    .Y(_0994_));
 sg13g2_nor3_1 _1905_ (.A(net708),
    .B(_0966_),
    .C(_0967_),
    .Y(_0995_));
 sg13g2_nor3_1 _1906_ (.A(net725),
    .B(_0993_),
    .C(_0994_),
    .Y(_0996_));
 sg13g2_nand3_1 _1907_ (.B(_0968_),
    .C(_0969_),
    .A(net727),
    .Y(_0997_));
 sg13g2_o21ai_1 _1908_ (.B1(net706),
    .Y(_0998_),
    .A1(_0995_),
    .A2(_0996_));
 sg13g2_nand3_1 _1909_ (.B(_0997_),
    .C(_0998_),
    .A(net704),
    .Y(_0999_));
 sg13g2_nand3_1 _1910_ (.B(_0970_),
    .C(_0971_),
    .A(net729),
    .Y(_1000_));
 sg13g2_nand3_1 _1911_ (.B(_0972_),
    .C(_0973_),
    .A(net731),
    .Y(_1001_));
 sg13g2_nand3_1 _1912_ (.B(_0999_),
    .C(_1000_),
    .A(net702),
    .Y(_1002_));
 sg13g2_nand3_1 _1913_ (.B(_1001_),
    .C(_1002_),
    .A(net699),
    .Y(_1003_));
 sg13g2_nand3_1 _1914_ (.B(_0988_),
    .C(_0989_),
    .A(net735),
    .Y(_1004_));
 sg13g2_o21ai_1 _1915_ (.B1(net713),
    .Y(_1005_),
    .A1(_0974_),
    .A2(_0975_));
 sg13g2_nand2b_1 _1916_ (.Y(_1006_),
    .B(net720),
    .A_N(\a[23] ));
 sg13g2_nand3_1 _1917_ (.B(_0976_),
    .C(_0977_),
    .A(net711),
    .Y(_1007_));
 sg13g2_nand3_1 _1918_ (.B(_1005_),
    .C(_1006_),
    .A(\ayayayayayaya.b[22] ),
    .Y(_1008_));
 sg13g2_nand3_1 _1919_ (.B(_1007_),
    .C(_1008_),
    .A(net722),
    .Y(_1009_));
 sg13g2_nand3_1 _1920_ (.B(_0978_),
    .C(_0979_),
    .A(net710),
    .Y(_1010_));
 sg13g2_nand3_1 _1921_ (.B(_0980_),
    .C(_0981_),
    .A(net708),
    .Y(_1011_));
 sg13g2_nand3_1 _1922_ (.B(_1009_),
    .C(_1010_),
    .A(net725),
    .Y(_1012_));
 sg13g2_nand3_1 _1923_ (.B(_1011_),
    .C(_1012_),
    .A(net727),
    .Y(_1013_));
 sg13g2_nand3_1 _1924_ (.B(_0982_),
    .C(_0983_),
    .A(net707),
    .Y(_1014_));
 sg13g2_nand3_1 _1925_ (.B(_0984_),
    .C(_0985_),
    .A(net704),
    .Y(_1015_));
 sg13g2_nand3_1 _1926_ (.B(_1013_),
    .C(_1014_),
    .A(net729),
    .Y(_1016_));
 sg13g2_nand3_1 _1927_ (.B(_1015_),
    .C(_1016_),
    .A(net732),
    .Y(_1017_));
 sg13g2_nand3_1 _1928_ (.B(_0986_),
    .C(_0987_),
    .A(net702),
    .Y(_1018_));
 sg13g2_nand3_1 _1929_ (.B(_0988_),
    .C(_0989_),
    .A(net699),
    .Y(_1019_));
 sg13g2_nand3_1 _1930_ (.B(_1017_),
    .C(_1018_),
    .A(net735),
    .Y(_1020_));
 sg13g2_nand3_1 _1931_ (.B(_1019_),
    .C(_1020_),
    .A(net738),
    .Y(_1021_));
 sg13g2_nand3_1 _1932_ (.B(_1003_),
    .C(_1004_),
    .A(net697),
    .Y(_1022_));
 sg13g2_nor2_1 _1933_ (.A(net712),
    .B(_0990_),
    .Y(_1023_));
 sg13g2_o21ai_1 _1934_ (.B1(_0762_),
    .Y(_1024_),
    .A1(net712),
    .A2(_0990_));
 sg13g2_o21ai_1 _1935_ (.B1(net723),
    .Y(_1025_),
    .A1(_0991_),
    .A2(_0992_));
 sg13g2_nor3_1 _1936_ (.A(net708),
    .B(_0993_),
    .C(_0994_),
    .Y(_1026_));
 sg13g2_a21oi_1 _1937_ (.A1(_1024_),
    .A2(_1025_),
    .Y(_1027_),
    .B1(net725));
 sg13g2_nor3_1 _1938_ (.A(net727),
    .B(_1026_),
    .C(_1027_),
    .Y(_1028_));
 sg13g2_nor3_1 _1939_ (.A(net706),
    .B(_0995_),
    .C(_0996_),
    .Y(_1029_));
 sg13g2_o21ai_1 _1940_ (.B1(net705),
    .Y(_1030_),
    .A1(_1028_),
    .A2(_1029_));
 sg13g2_nand3_1 _1941_ (.B(_0997_),
    .C(_0998_),
    .A(net729),
    .Y(_1031_));
 sg13g2_nand3_1 _1942_ (.B(_0999_),
    .C(_1000_),
    .A(net731),
    .Y(_1032_));
 sg13g2_nand3_1 _1943_ (.B(_1030_),
    .C(_1031_),
    .A(net702),
    .Y(_1033_));
 sg13g2_nand3_1 _1944_ (.B(_1032_),
    .C(_1033_),
    .A(net699),
    .Y(_1034_));
 sg13g2_nand3_1 _1945_ (.B(_1001_),
    .C(_1002_),
    .A(net735),
    .Y(_1035_));
 sg13g2_nand3_1 _1946_ (.B(_1003_),
    .C(_1004_),
    .A(net738),
    .Y(_1036_));
 sg13g2_nand3_1 _1947_ (.B(_1034_),
    .C(_1035_),
    .A(net697),
    .Y(_1037_));
 sg13g2_nand3_1 _1948_ (.B(_1036_),
    .C(_1037_),
    .A(net694),
    .Y(_1038_));
 sg13g2_nand3_1 _1949_ (.B(_1021_),
    .C(_1022_),
    .A(net743),
    .Y(_1039_));
 sg13g2_a21oi_1 _1950_ (.A1(_1005_),
    .A2(_1006_),
    .Y(_1040_),
    .B1(net721));
 sg13g2_nor2_1 _1951_ (.A(\a[22] ),
    .B(net711),
    .Y(_1041_));
 sg13g2_o21ai_1 _1952_ (.B1(net722),
    .Y(_1042_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_nand3_1 _1953_ (.B(_1007_),
    .C(_1008_),
    .A(net710),
    .Y(_1043_));
 sg13g2_nand3_1 _1954_ (.B(_1009_),
    .C(_1010_),
    .A(net708),
    .Y(_1044_));
 sg13g2_nand3_1 _1955_ (.B(_1042_),
    .C(_1043_),
    .A(net726),
    .Y(_1045_));
 sg13g2_nand3_1 _1956_ (.B(_1044_),
    .C(_1045_),
    .A(net728),
    .Y(_1046_));
 sg13g2_nand3_1 _1957_ (.B(_1011_),
    .C(_1012_),
    .A(net707),
    .Y(_1047_));
 sg13g2_nand3_1 _1958_ (.B(_1013_),
    .C(_1014_),
    .A(net705),
    .Y(_1048_));
 sg13g2_nand3_1 _1959_ (.B(_1046_),
    .C(_1047_),
    .A(net730),
    .Y(_1049_));
 sg13g2_nand3_1 _1960_ (.B(_1048_),
    .C(_1049_),
    .A(net732),
    .Y(_1050_));
 sg13g2_nand3_1 _1961_ (.B(_1015_),
    .C(_1016_),
    .A(net702),
    .Y(_1051_));
 sg13g2_nand3_1 _1962_ (.B(_1017_),
    .C(_1018_),
    .A(net700),
    .Y(_1052_));
 sg13g2_nand3_1 _1963_ (.B(_1050_),
    .C(_1051_),
    .A(net735),
    .Y(_1053_));
 sg13g2_nand2_1 _1964_ (.Y(_1054_),
    .A(_1052_),
    .B(_1053_));
 sg13g2_nand3_1 _1965_ (.B(_1052_),
    .C(_1053_),
    .A(net738),
    .Y(_1055_));
 sg13g2_nand3_1 _1966_ (.B(_1019_),
    .C(_1020_),
    .A(net697),
    .Y(_1056_));
 sg13g2_nand3_1 _1967_ (.B(_1021_),
    .C(_1022_),
    .A(net694),
    .Y(_1057_));
 sg13g2_nand3_1 _1968_ (.B(_1055_),
    .C(_1056_),
    .A(net742),
    .Y(_1058_));
 sg13g2_nand3_1 _1969_ (.B(_1057_),
    .C(_1058_),
    .A(net746),
    .Y(_1059_));
 sg13g2_nand3_1 _1970_ (.B(_1038_),
    .C(_1039_),
    .A(net689),
    .Y(_1060_));
 sg13g2_nand3_1 _1971_ (.B(net709),
    .C(_1023_),
    .A(net722),
    .Y(_1061_));
 sg13g2_nand3_1 _1972_ (.B(_1024_),
    .C(_1025_),
    .A(net725),
    .Y(_1062_));
 sg13g2_a21oi_1 _1973_ (.A1(_1061_),
    .A2(_1062_),
    .Y(_1063_),
    .B1(net728));
 sg13g2_nor3_1 _1974_ (.A(net707),
    .B(_1026_),
    .C(_1027_),
    .Y(_1064_));
 sg13g2_nor3_1 _1975_ (.A(net704),
    .B(_1028_),
    .C(_1029_),
    .Y(_1065_));
 sg13g2_nor3_1 _1976_ (.A(net729),
    .B(_1063_),
    .C(_1064_),
    .Y(_1066_));
 sg13g2_nand3_1 _1977_ (.B(_1030_),
    .C(_1031_),
    .A(net731),
    .Y(_1067_));
 sg13g2_o21ai_1 _1978_ (.B1(net702),
    .Y(_1068_),
    .A1(_1065_),
    .A2(_1066_));
 sg13g2_nand3_1 _1979_ (.B(_1067_),
    .C(_1068_),
    .A(net700),
    .Y(_1069_));
 sg13g2_nand3_1 _1980_ (.B(_1032_),
    .C(_1033_),
    .A(net735),
    .Y(_1070_));
 sg13g2_nand2_1 _1981_ (.Y(_1071_),
    .A(_1069_),
    .B(_1070_));
 sg13g2_nand3_1 _1982_ (.B(_1034_),
    .C(_1035_),
    .A(net738),
    .Y(_1072_));
 sg13g2_nand3_1 _1983_ (.B(_1069_),
    .C(_1070_),
    .A(_0813_),
    .Y(_1073_));
 sg13g2_nand3_1 _1984_ (.B(_1072_),
    .C(_1073_),
    .A(net693),
    .Y(_1074_));
 sg13g2_nand3_1 _1985_ (.B(_1036_),
    .C(_1037_),
    .A(net742),
    .Y(_1075_));
 sg13g2_nand3_1 _1986_ (.B(_1038_),
    .C(_1039_),
    .A(net746),
    .Y(_1076_));
 sg13g2_nand3_1 _1987_ (.B(_1074_),
    .C(_1075_),
    .A(net689),
    .Y(_1077_));
 sg13g2_nand3_1 _1988_ (.B(_1076_),
    .C(_1077_),
    .A(net686),
    .Y(_1078_));
 sg13g2_nand3_1 _1989_ (.B(_1059_),
    .C(_1060_),
    .A(net751),
    .Y(_1079_));
 sg13g2_o21ai_1 _1990_ (.B1(net710),
    .Y(_1080_),
    .A1(_1040_),
    .A2(_1041_));
 sg13g2_nand2b_1 _1991_ (.Y(_1081_),
    .B(net722),
    .A_N(\a[21] ));
 sg13g2_nand3_1 _1992_ (.B(_1042_),
    .C(_1043_),
    .A(net708),
    .Y(_1082_));
 sg13g2_nand3_1 _1993_ (.B(_1080_),
    .C(_1081_),
    .A(net726),
    .Y(_1083_));
 sg13g2_nand3_1 _1994_ (.B(_1082_),
    .C(_1083_),
    .A(net728),
    .Y(_1084_));
 sg13g2_nand3_1 _1995_ (.B(_1044_),
    .C(_1045_),
    .A(net707),
    .Y(_1085_));
 sg13g2_nand3_1 _1996_ (.B(_1046_),
    .C(_1047_),
    .A(net705),
    .Y(_1086_));
 sg13g2_nand3_1 _1997_ (.B(_1084_),
    .C(_1085_),
    .A(net730),
    .Y(_1087_));
 sg13g2_nand3_1 _1998_ (.B(_1086_),
    .C(_1087_),
    .A(net733),
    .Y(_1088_));
 sg13g2_nand3_1 _1999_ (.B(_1048_),
    .C(_1049_),
    .A(net703),
    .Y(_1089_));
 sg13g2_nand3_1 _2000_ (.B(_1050_),
    .C(_1051_),
    .A(net700),
    .Y(_1090_));
 sg13g2_nand3_1 _2001_ (.B(_1088_),
    .C(_1089_),
    .A(net736),
    .Y(_1091_));
 sg13g2_nand3_1 _2002_ (.B(_1090_),
    .C(_1091_),
    .A(net738),
    .Y(_1092_));
 sg13g2_nand3_1 _2003_ (.B(_1052_),
    .C(_1053_),
    .A(net697),
    .Y(_1093_));
 sg13g2_nand3_1 _2004_ (.B(_1055_),
    .C(_1056_),
    .A(net693),
    .Y(_1094_));
 sg13g2_nand3_1 _2005_ (.B(_1092_),
    .C(_1093_),
    .A(net742),
    .Y(_1095_));
 sg13g2_nand3_1 _2006_ (.B(_1094_),
    .C(_1095_),
    .A(net746),
    .Y(_1096_));
 sg13g2_nand3_1 _2007_ (.B(_1057_),
    .C(_1058_),
    .A(net689),
    .Y(_1097_));
 sg13g2_nand3_1 _2008_ (.B(_1059_),
    .C(_1060_),
    .A(net686),
    .Y(_1098_));
 sg13g2_nand3_1 _2009_ (.B(_1096_),
    .C(_1097_),
    .A(net750),
    .Y(_1099_));
 sg13g2_nand3_1 _2010_ (.B(_1098_),
    .C(_1099_),
    .A(net755),
    .Y(_1100_));
 sg13g2_nand3_1 _2011_ (.B(_1078_),
    .C(_1079_),
    .A(net682),
    .Y(_1101_));
 sg13g2_o21ai_1 _2012_ (.B1(\ayayayayayaya.b[18] ),
    .Y(_1102_),
    .A1(_1063_),
    .A2(_1064_));
 sg13g2_nand3_1 _2013_ (.B(net726),
    .C(_1023_),
    .A(net722),
    .Y(_1103_));
 sg13g2_nor2_1 _2014_ (.A(net727),
    .B(_1103_),
    .Y(_1104_));
 sg13g2_a21oi_1 _2015_ (.A1(_1061_),
    .A2(_1062_),
    .Y(_1105_),
    .B1(net706));
 sg13g2_o21ai_1 _2016_ (.B1(net704),
    .Y(_1106_),
    .A1(_1104_),
    .A2(_1105_));
 sg13g2_a21oi_1 _2017_ (.A1(_1102_),
    .A2(_1106_),
    .Y(_1107_),
    .B1(net731));
 sg13g2_nor3_1 _2018_ (.A(net702),
    .B(_1065_),
    .C(_1066_),
    .Y(_1108_));
 sg13g2_o21ai_1 _2019_ (.B1(net699),
    .Y(_1109_),
    .A1(_1107_),
    .A2(_1108_));
 sg13g2_nand3_1 _2020_ (.B(_1067_),
    .C(_1068_),
    .A(net735),
    .Y(_1110_));
 sg13g2_nand2_1 _2021_ (.Y(_1111_),
    .A(_1109_),
    .B(_1110_));
 sg13g2_nand3_1 _2022_ (.B(_1069_),
    .C(_1070_),
    .A(net739),
    .Y(_1112_));
 sg13g2_nand3_1 _2023_ (.B(_1109_),
    .C(_1110_),
    .A(net697),
    .Y(_1113_));
 sg13g2_nand3_1 _2024_ (.B(_1112_),
    .C(_1113_),
    .A(net693),
    .Y(_1114_));
 sg13g2_nand3_1 _2025_ (.B(_1072_),
    .C(_1073_),
    .A(net742),
    .Y(_1115_));
 sg13g2_nand3_1 _2026_ (.B(_1074_),
    .C(_1075_),
    .A(net746),
    .Y(_1116_));
 sg13g2_nand3_1 _2027_ (.B(_1114_),
    .C(_1115_),
    .A(net689),
    .Y(_1117_));
 sg13g2_nand3_1 _2028_ (.B(_1116_),
    .C(_1117_),
    .A(net686),
    .Y(_1118_));
 sg13g2_nand3_1 _2029_ (.B(_1076_),
    .C(_1077_),
    .A(net751),
    .Y(_1119_));
 sg13g2_nand3_1 _2030_ (.B(_1078_),
    .C(_1079_),
    .A(net755),
    .Y(_1120_));
 sg13g2_nand3_1 _2031_ (.B(_1118_),
    .C(_1119_),
    .A(net682),
    .Y(_1121_));
 sg13g2_nand3_1 _2032_ (.B(_1120_),
    .C(_1121_),
    .A(net679),
    .Y(_1122_));
 sg13g2_nand3_1 _2033_ (.B(_1100_),
    .C(_1101_),
    .A(net761),
    .Y(_1123_));
 sg13g2_a21oi_1 _2034_ (.A1(_1080_),
    .A2(_1081_),
    .Y(_1124_),
    .B1(net726));
 sg13g2_nor2_1 _2035_ (.A(\a[20] ),
    .B(net708),
    .Y(_1125_));
 sg13g2_o21ai_1 _2036_ (.B1(net728),
    .Y(_1126_),
    .A1(_1124_),
    .A2(_1125_));
 sg13g2_nand3_1 _2037_ (.B(_1082_),
    .C(_1083_),
    .A(net707),
    .Y(_1127_));
 sg13g2_nand3_1 _2038_ (.B(_1084_),
    .C(_1085_),
    .A(net705),
    .Y(_1128_));
 sg13g2_nand3_1 _2039_ (.B(_1126_),
    .C(_1127_),
    .A(net730),
    .Y(_1129_));
 sg13g2_nand3_1 _2040_ (.B(_1128_),
    .C(_1129_),
    .A(net733),
    .Y(_1130_));
 sg13g2_nand3_1 _2041_ (.B(_1086_),
    .C(_1087_),
    .A(net703),
    .Y(_1131_));
 sg13g2_nand3_1 _2042_ (.B(_1088_),
    .C(_1089_),
    .A(net700),
    .Y(_1132_));
 sg13g2_nand3_1 _2043_ (.B(_1130_),
    .C(_1131_),
    .A(net736),
    .Y(_1133_));
 sg13g2_nand3_1 _2044_ (.B(_1132_),
    .C(_1133_),
    .A(net740),
    .Y(_1134_));
 sg13g2_nand3_1 _2045_ (.B(_1090_),
    .C(_1091_),
    .A(net698),
    .Y(_1135_));
 sg13g2_nand3_1 _2046_ (.B(_1092_),
    .C(_1093_),
    .A(net693),
    .Y(_1136_));
 sg13g2_nand3_1 _2047_ (.B(_1134_),
    .C(_1135_),
    .A(net744),
    .Y(_1137_));
 sg13g2_nand3_1 _2048_ (.B(_1136_),
    .C(_1137_),
    .A(net746),
    .Y(_1138_));
 sg13g2_nand3_1 _2049_ (.B(_1094_),
    .C(_1095_),
    .A(net690),
    .Y(_1139_));
 sg13g2_nand3_1 _2050_ (.B(_1096_),
    .C(_1097_),
    .A(net687),
    .Y(_1140_));
 sg13g2_nand3_1 _2051_ (.B(_1138_),
    .C(_1139_),
    .A(net750),
    .Y(_1141_));
 sg13g2_nand3_1 _2052_ (.B(_1140_),
    .C(_1141_),
    .A(net756),
    .Y(_1142_));
 sg13g2_nand3_1 _2053_ (.B(_1098_),
    .C(_1099_),
    .A(net683),
    .Y(_1143_));
 sg13g2_nand3_1 _2054_ (.B(_1100_),
    .C(_1101_),
    .A(_0839_),
    .Y(_1144_));
 sg13g2_nand3_1 _2055_ (.B(_1142_),
    .C(_1143_),
    .A(net761),
    .Y(_1145_));
 sg13g2_nand3_1 _2056_ (.B(_1144_),
    .C(_1145_),
    .A(net766),
    .Y(_1146_));
 sg13g2_nand3_1 _2057_ (.B(_1122_),
    .C(_1123_),
    .A(net677),
    .Y(_1147_));
 sg13g2_nor2_1 _2058_ (.A(net706),
    .B(_1103_),
    .Y(_1148_));
 sg13g2_nand2_1 _2059_ (.Y(_1149_),
    .A(net704),
    .B(_1148_));
 sg13g2_o21ai_1 _2060_ (.B1(net729),
    .Y(_1150_),
    .A1(_1104_),
    .A2(_1105_));
 sg13g2_a21oi_1 _2061_ (.A1(_1149_),
    .A2(_1150_),
    .Y(_1151_),
    .B1(net731));
 sg13g2_a21oi_1 _2062_ (.A1(_1102_),
    .A2(_1106_),
    .Y(_1152_),
    .B1(net703));
 sg13g2_nor3_1 _2063_ (.A(net700),
    .B(_1107_),
    .C(_1108_),
    .Y(_1153_));
 sg13g2_nor3_1 _2064_ (.A(net736),
    .B(_1151_),
    .C(_1152_),
    .Y(_1154_));
 sg13g2_nand3_1 _2065_ (.B(_1109_),
    .C(_1110_),
    .A(net738),
    .Y(_1155_));
 sg13g2_o21ai_1 _2066_ (.B1(net697),
    .Y(_1156_),
    .A1(_1153_),
    .A2(_1154_));
 sg13g2_nand3_1 _2067_ (.B(_1155_),
    .C(_1156_),
    .A(net694),
    .Y(_1157_));
 sg13g2_nand3_1 _2068_ (.B(_1112_),
    .C(_1113_),
    .A(net742),
    .Y(_1158_));
 sg13g2_nand3_1 _2069_ (.B(_1114_),
    .C(_1115_),
    .A(net747),
    .Y(_1159_));
 sg13g2_nand3_1 _2070_ (.B(_1157_),
    .C(_1158_),
    .A(net689),
    .Y(_1160_));
 sg13g2_nand3_1 _2071_ (.B(_1159_),
    .C(_1160_),
    .A(net686),
    .Y(_1161_));
 sg13g2_nand3_1 _2072_ (.B(_1116_),
    .C(_1117_),
    .A(net750),
    .Y(_1162_));
 sg13g2_nand3_1 _2073_ (.B(_1118_),
    .C(_1119_),
    .A(net755),
    .Y(_1163_));
 sg13g2_nand3_1 _2074_ (.B(_1161_),
    .C(_1162_),
    .A(net682),
    .Y(_1164_));
 sg13g2_nand3_1 _2075_ (.B(_1163_),
    .C(_1164_),
    .A(net679),
    .Y(_1165_));
 sg13g2_nand3_1 _2076_ (.B(_1120_),
    .C(_1121_),
    .A(net760),
    .Y(_1166_));
 sg13g2_nand3_1 _2077_ (.B(_1122_),
    .C(_1123_),
    .A(net767),
    .Y(_1167_));
 sg13g2_nand3_1 _2078_ (.B(_1165_),
    .C(_1166_),
    .A(net676),
    .Y(_1168_));
 sg13g2_nand3_1 _2079_ (.B(_1167_),
    .C(_1168_),
    .A(net670),
    .Y(_1169_));
 sg13g2_nand3_1 _2080_ (.B(_1146_),
    .C(_1147_),
    .A(net771),
    .Y(_1170_));
 sg13g2_o21ai_1 _2081_ (.B1(net707),
    .Y(_1171_),
    .A1(_1124_),
    .A2(_1125_));
 sg13g2_nand2b_1 _2082_ (.Y(_1172_),
    .B(net728),
    .A_N(\a[19] ));
 sg13g2_nand3_1 _2083_ (.B(_1126_),
    .C(_1127_),
    .A(net705),
    .Y(_1173_));
 sg13g2_nand3_1 _2084_ (.B(_1171_),
    .C(_1172_),
    .A(net730),
    .Y(_1174_));
 sg13g2_nand3_1 _2085_ (.B(_1173_),
    .C(_1174_),
    .A(net733),
    .Y(_1175_));
 sg13g2_nand3_1 _2086_ (.B(_1128_),
    .C(_1129_),
    .A(net703),
    .Y(_1176_));
 sg13g2_nand3_1 _2087_ (.B(_1130_),
    .C(_1131_),
    .A(net701),
    .Y(_1177_));
 sg13g2_nand3_1 _2088_ (.B(_1175_),
    .C(_1176_),
    .A(net736),
    .Y(_1178_));
 sg13g2_nand3_1 _2089_ (.B(_1177_),
    .C(_1178_),
    .A(net740),
    .Y(_1179_));
 sg13g2_nand3_1 _2090_ (.B(_1132_),
    .C(_1133_),
    .A(net698),
    .Y(_1180_));
 sg13g2_nand3_1 _2091_ (.B(_1134_),
    .C(_1135_),
    .A(net695),
    .Y(_1181_));
 sg13g2_nand3_1 _2092_ (.B(_1179_),
    .C(_1180_),
    .A(net744),
    .Y(_1182_));
 sg13g2_nand3_1 _2093_ (.B(_1181_),
    .C(_1182_),
    .A(\ayayayayayaya.b[13] ),
    .Y(_1183_));
 sg13g2_nand3_1 _2094_ (.B(_1136_),
    .C(_1137_),
    .A(net690),
    .Y(_1184_));
 sg13g2_nand3_1 _2095_ (.B(_1138_),
    .C(_1139_),
    .A(net687),
    .Y(_1185_));
 sg13g2_nand3_1 _2096_ (.B(_1183_),
    .C(_1184_),
    .A(net750),
    .Y(_1186_));
 sg13g2_nand3_1 _2097_ (.B(_1185_),
    .C(_1186_),
    .A(net756),
    .Y(_1187_));
 sg13g2_nand3_1 _2098_ (.B(_1140_),
    .C(_1141_),
    .A(net683),
    .Y(_1188_));
 sg13g2_nand3_1 _2099_ (.B(_1142_),
    .C(_1143_),
    .A(_0839_),
    .Y(_1189_));
 sg13g2_nand3_1 _2100_ (.B(_1187_),
    .C(_1188_),
    .A(net761),
    .Y(_1190_));
 sg13g2_nand3_1 _2101_ (.B(_1189_),
    .C(_1190_),
    .A(net765),
    .Y(_1191_));
 sg13g2_nand3_1 _2102_ (.B(_1144_),
    .C(_1145_),
    .A(net678),
    .Y(_1192_));
 sg13g2_nand3_1 _2103_ (.B(_1146_),
    .C(_1147_),
    .A(net671),
    .Y(_1193_));
 sg13g2_nand3_1 _2104_ (.B(_1191_),
    .C(_1192_),
    .A(net771),
    .Y(_1194_));
 sg13g2_nand3_1 _2105_ (.B(_1193_),
    .C(_1194_),
    .A(net776),
    .Y(_1195_));
 sg13g2_nand3_1 _2106_ (.B(_1169_),
    .C(_1170_),
    .A(net667),
    .Y(_1196_));
 sg13g2_a21o_1 _2107_ (.A2(_1148_),
    .A1(\ayayayayayaya.b[18] ),
    .B1(net731),
    .X(_1197_));
 sg13g2_nand3_1 _2108_ (.B(_1149_),
    .C(_1150_),
    .A(net731),
    .Y(_1198_));
 sg13g2_nor3_1 _2109_ (.A(net700),
    .B(_1151_),
    .C(_1152_),
    .Y(_1199_));
 sg13g2_a21oi_1 _2110_ (.A1(_1197_),
    .A2(_1198_),
    .Y(_1200_),
    .B1(net735));
 sg13g2_nor2_1 _2111_ (.A(_1199_),
    .B(_1200_),
    .Y(_1201_));
 sg13g2_nor3_1 _2112_ (.A(net739),
    .B(_1199_),
    .C(_1200_),
    .Y(_1202_));
 sg13g2_nor3_1 _2113_ (.A(net698),
    .B(_1153_),
    .C(_1154_),
    .Y(_1203_));
 sg13g2_o21ai_1 _2114_ (.B1(net693),
    .Y(_1204_),
    .A1(_1202_),
    .A2(_1203_));
 sg13g2_nand3_1 _2115_ (.B(_1155_),
    .C(_1156_),
    .A(net742),
    .Y(_1205_));
 sg13g2_nand3_1 _2116_ (.B(_1157_),
    .C(_1158_),
    .A(net747),
    .Y(_1206_));
 sg13g2_nand3_1 _2117_ (.B(_1204_),
    .C(_1205_),
    .A(net690),
    .Y(_1207_));
 sg13g2_nand3_1 _2118_ (.B(_1206_),
    .C(_1207_),
    .A(net688),
    .Y(_1208_));
 sg13g2_nand3_1 _2119_ (.B(_1159_),
    .C(_1160_),
    .A(net750),
    .Y(_1209_));
 sg13g2_nand3_1 _2120_ (.B(_1161_),
    .C(_1162_),
    .A(net755),
    .Y(_1210_));
 sg13g2_nand3_1 _2121_ (.B(_1208_),
    .C(_1209_),
    .A(net683),
    .Y(_1211_));
 sg13g2_nand3_1 _2122_ (.B(_1210_),
    .C(_1211_),
    .A(net679),
    .Y(_1212_));
 sg13g2_nand3_1 _2123_ (.B(_1163_),
    .C(_1164_),
    .A(net760),
    .Y(_1213_));
 sg13g2_nand3_1 _2124_ (.B(_1165_),
    .C(_1166_),
    .A(net766),
    .Y(_1214_));
 sg13g2_nand3_1 _2125_ (.B(_1212_),
    .C(_1213_),
    .A(net676),
    .Y(_1215_));
 sg13g2_nand3_1 _2126_ (.B(_1214_),
    .C(_1215_),
    .A(net670),
    .Y(_1216_));
 sg13g2_nand3_1 _2127_ (.B(_1167_),
    .C(_1168_),
    .A(net771),
    .Y(_1217_));
 sg13g2_nand3_1 _2128_ (.B(_1169_),
    .C(_1170_),
    .A(net777),
    .Y(_1218_));
 sg13g2_nand3_1 _2129_ (.B(_1216_),
    .C(_1217_),
    .A(net667),
    .Y(_1219_));
 sg13g2_nand3_1 _2130_ (.B(_1218_),
    .C(_1219_),
    .A(net662),
    .Y(_1220_));
 sg13g2_nand3_1 _2131_ (.B(_1195_),
    .C(_1196_),
    .A(net783),
    .Y(_1221_));
 sg13g2_a21oi_1 _2132_ (.A1(_1171_),
    .A2(_1172_),
    .Y(_1222_),
    .B1(net730));
 sg13g2_nor2_1 _2133_ (.A(\a[18] ),
    .B(net705),
    .Y(_1223_));
 sg13g2_o21ai_1 _2134_ (.B1(net733),
    .Y(_1224_),
    .A1(_1222_),
    .A2(_1223_));
 sg13g2_nand3_1 _2135_ (.B(_1173_),
    .C(_1174_),
    .A(net703),
    .Y(_1225_));
 sg13g2_nand3_1 _2136_ (.B(_1175_),
    .C(_1176_),
    .A(net701),
    .Y(_1226_));
 sg13g2_nand3_1 _2137_ (.B(_1224_),
    .C(_1225_),
    .A(net736),
    .Y(_1227_));
 sg13g2_nand3_1 _2138_ (.B(_1226_),
    .C(_1227_),
    .A(net740),
    .Y(_1228_));
 sg13g2_nand3_1 _2139_ (.B(_1177_),
    .C(_1178_),
    .A(net698),
    .Y(_1229_));
 sg13g2_nand3_1 _2140_ (.B(_1179_),
    .C(_1180_),
    .A(net695),
    .Y(_1230_));
 sg13g2_nand3_1 _2141_ (.B(_1228_),
    .C(_1229_),
    .A(net744),
    .Y(_1231_));
 sg13g2_nand3_1 _2142_ (.B(_1230_),
    .C(_1231_),
    .A(\ayayayayayaya.b[13] ),
    .Y(_1232_));
 sg13g2_nand3_1 _2143_ (.B(_1181_),
    .C(_1182_),
    .A(net691),
    .Y(_1233_));
 sg13g2_nand3_1 _2144_ (.B(_1183_),
    .C(_1184_),
    .A(net687),
    .Y(_1234_));
 sg13g2_nand3_1 _2145_ (.B(_1232_),
    .C(_1233_),
    .A(net752),
    .Y(_1235_));
 sg13g2_nand3_1 _2146_ (.B(_1234_),
    .C(_1235_),
    .A(net756),
    .Y(_1236_));
 sg13g2_nand3_1 _2147_ (.B(_1185_),
    .C(_1186_),
    .A(net683),
    .Y(_1237_));
 sg13g2_nand3_1 _2148_ (.B(_1187_),
    .C(_1188_),
    .A(net680),
    .Y(_1238_));
 sg13g2_nand3_1 _2149_ (.B(_1236_),
    .C(_1237_),
    .A(net760),
    .Y(_1239_));
 sg13g2_nand3_1 _2150_ (.B(_1238_),
    .C(_1239_),
    .A(net765),
    .Y(_1240_));
 sg13g2_nand3_1 _2151_ (.B(_1189_),
    .C(_1190_),
    .A(net678),
    .Y(_1241_));
 sg13g2_nand3_1 _2152_ (.B(_1191_),
    .C(_1192_),
    .A(net671),
    .Y(_1242_));
 sg13g2_nand3_1 _2153_ (.B(_1240_),
    .C(_1241_),
    .A(net770),
    .Y(_1243_));
 sg13g2_nand3_1 _2154_ (.B(_1242_),
    .C(_1243_),
    .A(net777),
    .Y(_1244_));
 sg13g2_nand3_1 _2155_ (.B(_1193_),
    .C(_1194_),
    .A(net666),
    .Y(_1245_));
 sg13g2_nand3_1 _2156_ (.B(_1195_),
    .C(_1196_),
    .A(net661),
    .Y(_1246_));
 sg13g2_nand3_1 _2157_ (.B(_1244_),
    .C(_1245_),
    .A(net782),
    .Y(_1247_));
 sg13g2_nand3_1 _2158_ (.B(_1246_),
    .C(_1247_),
    .A(net791),
    .Y(_1248_));
 sg13g2_nand3_1 _2159_ (.B(_1220_),
    .C(_1221_),
    .A(net657),
    .Y(_1249_));
 sg13g2_nand3_1 _2160_ (.B(net731),
    .C(_1148_),
    .A(\ayayayayayaya.b[18] ),
    .Y(_1250_));
 sg13g2_and2_1 _2161_ (.A(net699),
    .B(_1250_),
    .X(_1251_));
 sg13g2_a21oi_1 _2162_ (.A1(_1197_),
    .A2(_1198_),
    .Y(_1252_),
    .B1(net699));
 sg13g2_nor2_1 _2163_ (.A(_1251_),
    .B(_1252_),
    .Y(_1253_));
 sg13g2_nor3_1 _2164_ (.A(net738),
    .B(_1251_),
    .C(_1252_),
    .Y(_1254_));
 sg13g2_nor3_1 _2165_ (.A(net698),
    .B(_1199_),
    .C(_1200_),
    .Y(_1255_));
 sg13g2_nor3_1 _2166_ (.A(net694),
    .B(_1202_),
    .C(_1203_),
    .Y(_1256_));
 sg13g2_nor3_1 _2167_ (.A(net743),
    .B(_1254_),
    .C(_1255_),
    .Y(_1257_));
 sg13g2_nand3_1 _2168_ (.B(_1204_),
    .C(_1205_),
    .A(net746),
    .Y(_1258_));
 sg13g2_o21ai_1 _2169_ (.B1(net689),
    .Y(_1259_),
    .A1(_1256_),
    .A2(_1257_));
 sg13g2_nand3_1 _2170_ (.B(_1258_),
    .C(_1259_),
    .A(net686),
    .Y(_1260_));
 sg13g2_nand3_1 _2171_ (.B(_1206_),
    .C(_1207_),
    .A(net751),
    .Y(_1261_));
 sg13g2_nand3_1 _2172_ (.B(_1208_),
    .C(_1209_),
    .A(net755),
    .Y(_1262_));
 sg13g2_nand3_1 _2173_ (.B(_1260_),
    .C(_1261_),
    .A(net682),
    .Y(_1263_));
 sg13g2_nand3_1 _2174_ (.B(_1262_),
    .C(_1263_),
    .A(net679),
    .Y(_1264_));
 sg13g2_nand3_1 _2175_ (.B(_1210_),
    .C(_1211_),
    .A(net760),
    .Y(_1265_));
 sg13g2_nand3_1 _2176_ (.B(_1212_),
    .C(_1213_),
    .A(net765),
    .Y(_1266_));
 sg13g2_nand3_1 _2177_ (.B(_1264_),
    .C(_1265_),
    .A(net676),
    .Y(_1267_));
 sg13g2_nand3_1 _2178_ (.B(_1266_),
    .C(_1267_),
    .A(net670),
    .Y(_1268_));
 sg13g2_nand3_1 _2179_ (.B(_1214_),
    .C(_1215_),
    .A(net771),
    .Y(_1269_));
 sg13g2_nand3_1 _2180_ (.B(_1216_),
    .C(_1217_),
    .A(net777),
    .Y(_1270_));
 sg13g2_nand3_1 _2181_ (.B(_1268_),
    .C(_1269_),
    .A(net667),
    .Y(_1271_));
 sg13g2_nand3_1 _2182_ (.B(_1270_),
    .C(_1271_),
    .A(net662),
    .Y(_1272_));
 sg13g2_nand3_1 _2183_ (.B(_1218_),
    .C(_1219_),
    .A(net783),
    .Y(_1273_));
 sg13g2_nand3_1 _2184_ (.B(_1220_),
    .C(_1221_),
    .A(net791),
    .Y(_1274_));
 sg13g2_nand3_1 _2185_ (.B(_1272_),
    .C(_1273_),
    .A(net657),
    .Y(_1275_));
 sg13g2_nand3_1 _2186_ (.B(_1274_),
    .C(_1275_),
    .A(net651),
    .Y(_1276_));
 sg13g2_nand3_1 _2187_ (.B(_1248_),
    .C(_1249_),
    .A(net797),
    .Y(_1277_));
 sg13g2_o21ai_1 _2188_ (.B1(net703),
    .Y(_1278_),
    .A1(_1222_),
    .A2(_1223_));
 sg13g2_nand2b_1 _2189_ (.Y(_1279_),
    .B(net734),
    .A_N(\a[17] ));
 sg13g2_nand3_1 _2190_ (.B(_1224_),
    .C(_1225_),
    .A(net701),
    .Y(_1280_));
 sg13g2_nand3_1 _2191_ (.B(_1278_),
    .C(_1279_),
    .A(net737),
    .Y(_1281_));
 sg13g2_nand3_1 _2192_ (.B(_1280_),
    .C(_1281_),
    .A(net740),
    .Y(_1282_));
 sg13g2_nand3_1 _2193_ (.B(_1226_),
    .C(_1227_),
    .A(net698),
    .Y(_1283_));
 sg13g2_nand3_1 _2194_ (.B(_1228_),
    .C(_1229_),
    .A(net695),
    .Y(_1284_));
 sg13g2_nand3_1 _2195_ (.B(_1282_),
    .C(_1283_),
    .A(net745),
    .Y(_1285_));
 sg13g2_nand3_1 _2196_ (.B(_1284_),
    .C(_1285_),
    .A(net748),
    .Y(_1286_));
 sg13g2_nand3_1 _2197_ (.B(_1230_),
    .C(_1231_),
    .A(net691),
    .Y(_1287_));
 sg13g2_nand3_1 _2198_ (.B(_1232_),
    .C(_1233_),
    .A(net687),
    .Y(_1288_));
 sg13g2_nand3_1 _2199_ (.B(_1286_),
    .C(_1287_),
    .A(net752),
    .Y(_1289_));
 sg13g2_nand3_1 _2200_ (.B(_1288_),
    .C(_1289_),
    .A(net756),
    .Y(_1290_));
 sg13g2_nand3_1 _2201_ (.B(_1234_),
    .C(_1235_),
    .A(net684),
    .Y(_1291_));
 sg13g2_nand3_1 _2202_ (.B(_1236_),
    .C(_1237_),
    .A(net680),
    .Y(_1292_));
 sg13g2_nand3_1 _2203_ (.B(_1290_),
    .C(_1291_),
    .A(net761),
    .Y(_1293_));
 sg13g2_nand3_1 _2204_ (.B(_1292_),
    .C(_1293_),
    .A(net766),
    .Y(_1294_));
 sg13g2_nand3_1 _2205_ (.B(_1238_),
    .C(_1239_),
    .A(net676),
    .Y(_1295_));
 sg13g2_nand3_1 _2206_ (.B(_1240_),
    .C(_1241_),
    .A(net670),
    .Y(_1296_));
 sg13g2_nand3_1 _2207_ (.B(_1294_),
    .C(_1295_),
    .A(net770),
    .Y(_1297_));
 sg13g2_nand3_1 _2208_ (.B(_1296_),
    .C(_1297_),
    .A(net777),
    .Y(_1298_));
 sg13g2_nand3_1 _2209_ (.B(_1242_),
    .C(_1243_),
    .A(net666),
    .Y(_1299_));
 sg13g2_nand3_1 _2210_ (.B(_1244_),
    .C(_1245_),
    .A(net662),
    .Y(_1300_));
 sg13g2_nand3_1 _2211_ (.B(_1298_),
    .C(_1299_),
    .A(net783),
    .Y(_1301_));
 sg13g2_nand3_1 _2212_ (.B(_1300_),
    .C(_1301_),
    .A(net790),
    .Y(_1302_));
 sg13g2_nand3_1 _2213_ (.B(_1246_),
    .C(_1247_),
    .A(net657),
    .Y(_1303_));
 sg13g2_nand3_1 _2214_ (.B(_1248_),
    .C(_1249_),
    .A(net651),
    .Y(_1304_));
 sg13g2_nand3_1 _2215_ (.B(_1302_),
    .C(_1303_),
    .A(net797),
    .Y(_1305_));
 sg13g2_nand3_1 _2216_ (.B(_1304_),
    .C(_1305_),
    .A(net804),
    .Y(_1306_));
 sg13g2_nand3_1 _2217_ (.B(_1276_),
    .C(_1277_),
    .A(net644),
    .Y(_1307_));
 sg13g2_nor2_2 _2218_ (.A(net700),
    .B(_1250_),
    .Y(_1308_));
 sg13g2_o21ai_1 _2219_ (.B1(net697),
    .Y(_1309_),
    .A1(net699),
    .A2(_1250_));
 sg13g2_o21ai_1 _2220_ (.B1(net738),
    .Y(_1310_),
    .A1(_1251_),
    .A2(_1252_));
 sg13g2_nor3_1 _2221_ (.A(net693),
    .B(_1254_),
    .C(_1255_),
    .Y(_1311_));
 sg13g2_a21oi_1 _2222_ (.A1(_1309_),
    .A2(_1310_),
    .Y(_1312_),
    .B1(net742));
 sg13g2_nor3_1 _2223_ (.A(net746),
    .B(_1311_),
    .C(_1312_),
    .Y(_1313_));
 sg13g2_nor3_1 _2224_ (.A(net689),
    .B(_1256_),
    .C(_1257_),
    .Y(_1314_));
 sg13g2_o21ai_1 _2225_ (.B1(net686),
    .Y(_1315_),
    .A1(_1313_),
    .A2(_1314_));
 sg13g2_nand3_1 _2226_ (.B(_1258_),
    .C(_1259_),
    .A(net751),
    .Y(_1316_));
 sg13g2_nand3_1 _2227_ (.B(_1260_),
    .C(_1261_),
    .A(net755),
    .Y(_1317_));
 sg13g2_nand3_1 _2228_ (.B(_1315_),
    .C(_1316_),
    .A(net682),
    .Y(_1318_));
 sg13g2_nand3_1 _2229_ (.B(_1317_),
    .C(_1318_),
    .A(net679),
    .Y(_1319_));
 sg13g2_nand3_1 _2230_ (.B(_1262_),
    .C(_1263_),
    .A(net760),
    .Y(_1320_));
 sg13g2_nand3_1 _2231_ (.B(_1264_),
    .C(_1265_),
    .A(net765),
    .Y(_1321_));
 sg13g2_nand3_1 _2232_ (.B(_1319_),
    .C(_1320_),
    .A(net676),
    .Y(_1322_));
 sg13g2_nand3_1 _2233_ (.B(_1321_),
    .C(_1322_),
    .A(net670),
    .Y(_1323_));
 sg13g2_nand3_1 _2234_ (.B(_1266_),
    .C(_1267_),
    .A(net770),
    .Y(_1324_));
 sg13g2_nand3_1 _2235_ (.B(_1268_),
    .C(_1269_),
    .A(net776),
    .Y(_1325_));
 sg13g2_nand3_1 _2236_ (.B(_1323_),
    .C(_1324_),
    .A(net666),
    .Y(_1326_));
 sg13g2_nand3_1 _2237_ (.B(_1325_),
    .C(_1326_),
    .A(net661),
    .Y(_1327_));
 sg13g2_nand3_1 _2238_ (.B(_1270_),
    .C(_1271_),
    .A(net783),
    .Y(_1328_));
 sg13g2_nand3_1 _2239_ (.B(_1272_),
    .C(_1273_),
    .A(net791),
    .Y(_1329_));
 sg13g2_nand3_1 _2240_ (.B(_1327_),
    .C(_1328_),
    .A(net657),
    .Y(_1330_));
 sg13g2_nand3_1 _2241_ (.B(_1329_),
    .C(_1330_),
    .A(net653),
    .Y(_1331_));
 sg13g2_nand3_1 _2242_ (.B(_1274_),
    .C(_1275_),
    .A(net797),
    .Y(_1332_));
 sg13g2_nand3_1 _2243_ (.B(_1276_),
    .C(_1277_),
    .A(net804),
    .Y(_1333_));
 sg13g2_nand3_1 _2244_ (.B(_1331_),
    .C(_1332_),
    .A(net644),
    .Y(_1334_));
 sg13g2_nand3_1 _2245_ (.B(_1333_),
    .C(_1334_),
    .A(net638),
    .Y(_1335_));
 sg13g2_nand3_1 _2246_ (.B(_1306_),
    .C(_1307_),
    .A(net810),
    .Y(_1336_));
 sg13g2_a21oi_1 _2247_ (.A1(_1278_),
    .A2(_1279_),
    .Y(_1337_),
    .B1(net737));
 sg13g2_nor2_1 _2248_ (.A(net831),
    .B(net701),
    .Y(_1338_));
 sg13g2_o21ai_1 _2249_ (.B1(net741),
    .Y(_1339_),
    .A1(_1337_),
    .A2(_1338_));
 sg13g2_nand3_1 _2250_ (.B(_1280_),
    .C(_1281_),
    .A(net698),
    .Y(_1340_));
 sg13g2_nand3_1 _2251_ (.B(_1282_),
    .C(_1283_),
    .A(net696),
    .Y(_1341_));
 sg13g2_nand3_1 _2252_ (.B(_1339_),
    .C(_1340_),
    .A(net745),
    .Y(_1342_));
 sg13g2_nand3_1 _2253_ (.B(_1341_),
    .C(_1342_),
    .A(net748),
    .Y(_1343_));
 sg13g2_nand3_1 _2254_ (.B(_1284_),
    .C(_1285_),
    .A(net692),
    .Y(_1344_));
 sg13g2_nand3_1 _2255_ (.B(_1286_),
    .C(_1287_),
    .A(net687),
    .Y(_1345_));
 sg13g2_nand3_1 _2256_ (.B(_1343_),
    .C(_1344_),
    .A(net749),
    .Y(_1346_));
 sg13g2_nand3_1 _2257_ (.B(_1345_),
    .C(_1346_),
    .A(net754),
    .Y(_1347_));
 sg13g2_nand3_1 _2258_ (.B(_1288_),
    .C(_1289_),
    .A(net684),
    .Y(_1348_));
 sg13g2_nand3_1 _2259_ (.B(_1290_),
    .C(_1291_),
    .A(net680),
    .Y(_1349_));
 sg13g2_nand3_1 _2260_ (.B(_1347_),
    .C(_1348_),
    .A(net761),
    .Y(_1350_));
 sg13g2_nand3_1 _2261_ (.B(_1349_),
    .C(_1350_),
    .A(net766),
    .Y(_1351_));
 sg13g2_nand3_1 _2262_ (.B(_1292_),
    .C(_1293_),
    .A(net677),
    .Y(_1352_));
 sg13g2_nand3_1 _2263_ (.B(_1294_),
    .C(_1295_),
    .A(net671),
    .Y(_1353_));
 sg13g2_nand3_1 _2264_ (.B(_1351_),
    .C(_1352_),
    .A(net772),
    .Y(_1354_));
 sg13g2_nand3_1 _2265_ (.B(_1353_),
    .C(_1354_),
    .A(net776),
    .Y(_1355_));
 sg13g2_nand3_1 _2266_ (.B(_1296_),
    .C(_1297_),
    .A(net667),
    .Y(_1356_));
 sg13g2_nand3_1 _2267_ (.B(_1298_),
    .C(_1299_),
    .A(net662),
    .Y(_1357_));
 sg13g2_nand3_1 _2268_ (.B(_1355_),
    .C(_1356_),
    .A(net782),
    .Y(_1358_));
 sg13g2_nand3_1 _2269_ (.B(_1357_),
    .C(_1358_),
    .A(net791),
    .Y(_1359_));
 sg13g2_nand3_1 _2270_ (.B(_1300_),
    .C(_1301_),
    .A(net657),
    .Y(_1360_));
 sg13g2_nand3_1 _2271_ (.B(_1302_),
    .C(_1303_),
    .A(net651),
    .Y(_1361_));
 sg13g2_nand3_1 _2272_ (.B(_1359_),
    .C(_1360_),
    .A(net796),
    .Y(_1362_));
 sg13g2_nand3_1 _2273_ (.B(_1361_),
    .C(_1362_),
    .A(net805),
    .Y(_1363_));
 sg13g2_nand3_1 _2274_ (.B(_1304_),
    .C(_1305_),
    .A(net643),
    .Y(_1364_));
 sg13g2_nand3_1 _2275_ (.B(_1306_),
    .C(_1307_),
    .A(net637),
    .Y(_1365_));
 sg13g2_nand3_1 _2276_ (.B(_1363_),
    .C(_1364_),
    .A(net811),
    .Y(_1366_));
 sg13g2_nand3_1 _2277_ (.B(_1365_),
    .C(_1366_),
    .A(net819),
    .Y(_1367_));
 sg13g2_nand3_1 _2278_ (.B(_1335_),
    .C(_1336_),
    .A(net631),
    .Y(_1368_));
 sg13g2_nand3_1 _2279_ (.B(_1367_),
    .C(_1368_),
    .A(net600),
    .Y(_1369_));
 sg13g2_nor2_1 _2280_ (.A(net822),
    .B(_0871_),
    .Y(_1370_));
 sg13g2_inv_1 _2281_ (.Y(_1371_),
    .A(net596));
 sg13g2_a21oi_1 _2282_ (.A1(net739),
    .A2(_1308_),
    .Y(_1372_),
    .B1(net742));
 sg13g2_a21oi_1 _2283_ (.A1(_1309_),
    .A2(_1310_),
    .Y(_1373_),
    .B1(net693));
 sg13g2_nor3_1 _2284_ (.A(net746),
    .B(_1372_),
    .C(_1373_),
    .Y(_1374_));
 sg13g2_nor3_1 _2285_ (.A(net690),
    .B(_1311_),
    .C(_1312_),
    .Y(_1375_));
 sg13g2_nor3_1 _2286_ (.A(net686),
    .B(_1313_),
    .C(_1314_),
    .Y(_1376_));
 sg13g2_nor3_1 _2287_ (.A(net750),
    .B(_1374_),
    .C(_1375_),
    .Y(_1377_));
 sg13g2_nand3_1 _2288_ (.B(_1315_),
    .C(_1316_),
    .A(net755),
    .Y(_1378_));
 sg13g2_o21ai_1 _2289_ (.B1(net682),
    .Y(_1379_),
    .A1(_1376_),
    .A2(_1377_));
 sg13g2_nand3_1 _2290_ (.B(_1378_),
    .C(_1379_),
    .A(net679),
    .Y(_1380_));
 sg13g2_nand3_1 _2291_ (.B(_1317_),
    .C(_1318_),
    .A(net760),
    .Y(_1381_));
 sg13g2_nand3_1 _2292_ (.B(_1319_),
    .C(_1320_),
    .A(net765),
    .Y(_1382_));
 sg13g2_nand3_1 _2293_ (.B(_1380_),
    .C(_1381_),
    .A(net676),
    .Y(_1383_));
 sg13g2_nand3_1 _2294_ (.B(_1382_),
    .C(_1383_),
    .A(net670),
    .Y(_1384_));
 sg13g2_nand3_1 _2295_ (.B(_1321_),
    .C(_1322_),
    .A(net770),
    .Y(_1385_));
 sg13g2_nand3_1 _2296_ (.B(_1323_),
    .C(_1324_),
    .A(net776),
    .Y(_1386_));
 sg13g2_nand3_1 _2297_ (.B(_1384_),
    .C(_1385_),
    .A(net666),
    .Y(_1387_));
 sg13g2_nand3_1 _2298_ (.B(_1386_),
    .C(_1387_),
    .A(net661),
    .Y(_1388_));
 sg13g2_nand3_1 _2299_ (.B(_1325_),
    .C(_1326_),
    .A(net782),
    .Y(_1389_));
 sg13g2_nand3_1 _2300_ (.B(_1327_),
    .C(_1328_),
    .A(net791),
    .Y(_1390_));
 sg13g2_nand3_1 _2301_ (.B(_1388_),
    .C(_1389_),
    .A(net656),
    .Y(_1391_));
 sg13g2_nand3_1 _2302_ (.B(_1390_),
    .C(_1391_),
    .A(net651),
    .Y(_1392_));
 sg13g2_nand3_1 _2303_ (.B(_1329_),
    .C(_1330_),
    .A(net797),
    .Y(_1393_));
 sg13g2_nand3_1 _2304_ (.B(_1331_),
    .C(_1332_),
    .A(net805),
    .Y(_1394_));
 sg13g2_nand3_1 _2305_ (.B(_1392_),
    .C(_1393_),
    .A(net644),
    .Y(_1395_));
 sg13g2_nand3_1 _2306_ (.B(_1394_),
    .C(_1395_),
    .A(net638),
    .Y(_1396_));
 sg13g2_nand3_1 _2307_ (.B(_1333_),
    .C(_1334_),
    .A(net810),
    .Y(_1397_));
 sg13g2_nand3_1 _2308_ (.B(_1335_),
    .C(_1336_),
    .A(net819),
    .Y(_1398_));
 sg13g2_nand3_1 _2309_ (.B(_1396_),
    .C(_1397_),
    .A(net631),
    .Y(_1399_));
 sg13g2_nand3_1 _2310_ (.B(_1398_),
    .C(_1399_),
    .A(net595),
    .Y(_1400_));
 sg13g2_nor2b_2 _2311_ (.A(net840),
    .B_N(net1),
    .Y(_1401_));
 sg13g2_and2_1 _2312_ (.A(_0869_),
    .B(_1401_),
    .X(_1402_));
 sg13g2_nor2_1 _2313_ (.A(net840),
    .B(net1),
    .Y(_1403_));
 sg13g2_and2_1 _2314_ (.A(_0869_),
    .B(_1403_),
    .X(_1404_));
 sg13g2_a22oi_1 _2315_ (.Y(_1405_),
    .B1(net619),
    .B2(net773),
    .A2(net623),
    .A1(net718));
 sg13g2_nor2_2 _2316_ (.A(net2),
    .B(net3),
    .Y(_1406_));
 sg13g2_or2_1 _2317_ (.X(_1407_),
    .B(net3),
    .A(net2));
 sg13g2_and2_1 _2318_ (.A(_1401_),
    .B(net838),
    .X(_1408_));
 sg13g2_nand2_2 _2319_ (.Y(_1409_),
    .A(_1401_),
    .B(net838));
 sg13g2_and2_1 _2320_ (.A(_1403_),
    .B(net838),
    .X(_1410_));
 sg13g2_nand2_1 _2321_ (.Y(_1411_),
    .A(_1403_),
    .B(net838));
 sg13g2_and2_1 _2322_ (.A(net841),
    .B(net838),
    .X(_1412_));
 sg13g2_and2_1 _2323_ (.A(\a[17] ),
    .B(net605),
    .X(_1413_));
 sg13g2_o21ai_1 _2324_ (.B1(net831),
    .Y(_1414_),
    .A1(net610),
    .A2(_1413_));
 sg13g2_nand3_1 _2325_ (.B(net831),
    .C(\a[17] ),
    .A(net842),
    .Y(_1415_));
 sg13g2_nor2b_2 _2326_ (.A(net3),
    .B_N(net2),
    .Y(_1416_));
 sg13g2_nand2b_2 _2327_ (.Y(_1417_),
    .B(net2),
    .A_N(net3));
 sg13g2_or2_1 _2328_ (.X(_1418_),
    .B(\a[17] ),
    .A(net830));
 sg13g2_nand3_1 _2329_ (.B(_1416_),
    .C(_1418_),
    .A(_1415_),
    .Y(_1419_));
 sg13g2_a21oi_1 _2330_ (.A1(net737),
    .A2(net615),
    .Y(_1420_),
    .B1(net848));
 sg13g2_nand4_1 _2331_ (.B(_1414_),
    .C(_1419_),
    .A(_1405_),
    .Y(_1421_),
    .D(_1420_));
 sg13g2_nor2b_2 _2332_ (.A(net1),
    .B_N(net840),
    .Y(_1422_));
 sg13g2_and2_1 _2333_ (.A(_0869_),
    .B(_1422_),
    .X(_1423_));
 sg13g2_nand2_1 _2334_ (.Y(_1424_),
    .A(_0869_),
    .B(_1422_));
 sg13g2_nor3_1 _2335_ (.A(_1337_),
    .B(_1338_),
    .C(net603),
    .Y(_1425_));
 sg13g2_nor2_1 _2336_ (.A(_1421_),
    .B(_1425_),
    .Y(_1426_));
 sg13g2_nand3_1 _2337_ (.B(_1400_),
    .C(_1426_),
    .A(_1369_),
    .Y(_1427_));
 sg13g2_and4_1 _2338_ (.A(net741),
    .B(net745),
    .C(net748),
    .D(_1308_),
    .X(_1428_));
 sg13g2_and3_1 _2339_ (.X(_1429_),
    .A(net752),
    .B(net684),
    .C(_1428_));
 sg13g2_nand2_1 _2340_ (.Y(_1430_),
    .A(net687),
    .B(_1428_));
 sg13g2_and4_1 _2341_ (.A(net740),
    .B(net744),
    .C(net691),
    .D(_1308_),
    .X(_1431_));
 sg13g2_nor3_1 _2342_ (.A(net690),
    .B(_1372_),
    .C(_1373_),
    .Y(_1432_));
 sg13g2_o21ai_1 _2343_ (.B1(net752),
    .Y(_1433_),
    .A1(_1431_),
    .A2(_1432_));
 sg13g2_a21oi_1 _2344_ (.A1(_1430_),
    .A2(_1433_),
    .Y(_1434_),
    .B1(net684));
 sg13g2_o21ai_1 _2345_ (.B1(net750),
    .Y(_1435_),
    .A1(_1374_),
    .A2(_1375_));
 sg13g2_o21ai_1 _2346_ (.B1(net687),
    .Y(_1436_),
    .A1(_1431_),
    .A2(_1432_));
 sg13g2_a21oi_1 _2347_ (.A1(_1430_),
    .A2(_1433_),
    .Y(_1437_),
    .B1(net756));
 sg13g2_a21oi_1 _2348_ (.A1(_1435_),
    .A2(_1436_),
    .Y(_1438_),
    .B1(net684));
 sg13g2_nor3_1 _2349_ (.A(net680),
    .B(_1437_),
    .C(_1438_),
    .Y(_1439_));
 sg13g2_nor3_1 _2350_ (.A(net761),
    .B(_1429_),
    .C(_1434_),
    .Y(_1440_));
 sg13g2_nand3_1 _2351_ (.B(net756),
    .C(_1428_),
    .A(net752),
    .Y(_1441_));
 sg13g2_and2_1 _2352_ (.A(net680),
    .B(_1441_),
    .X(_1442_));
 sg13g2_nor3_1 _2353_ (.A(net680),
    .B(_1429_),
    .C(_1434_),
    .Y(_1443_));
 sg13g2_nor3_1 _2354_ (.A(net766),
    .B(_1442_),
    .C(_1443_),
    .Y(_1444_));
 sg13g2_nor3_1 _2355_ (.A(net677),
    .B(_1439_),
    .C(_1440_),
    .Y(_1445_));
 sg13g2_a21oi_1 _2356_ (.A1(_1435_),
    .A2(_1436_),
    .Y(_1446_),
    .B1(net756));
 sg13g2_nor3_1 _2357_ (.A(net682),
    .B(_1376_),
    .C(_1377_),
    .Y(_1447_));
 sg13g2_o21ai_1 _2358_ (.B1(net679),
    .Y(_1448_),
    .A1(_1446_),
    .A2(_1447_));
 sg13g2_nand3_1 _2359_ (.B(_1378_),
    .C(_1379_),
    .A(net760),
    .Y(_1449_));
 sg13g2_nor2_1 _2360_ (.A(net681),
    .B(_1441_),
    .Y(_1450_));
 sg13g2_o21ai_1 _2361_ (.B1(net677),
    .Y(_1451_),
    .A1(net681),
    .A2(_1441_));
 sg13g2_o21ai_1 _2362_ (.B1(net766),
    .Y(_1452_),
    .A1(_1442_),
    .A2(_1443_));
 sg13g2_nor3_1 _2363_ (.A(net672),
    .B(_1444_),
    .C(_1445_),
    .Y(_1453_));
 sg13g2_a21oi_1 _2364_ (.A1(_1451_),
    .A2(_1452_),
    .Y(_1454_),
    .B1(net772));
 sg13g2_nor3_1 _2365_ (.A(net778),
    .B(_1453_),
    .C(_1454_),
    .Y(_1455_));
 sg13g2_nor3_1 _2366_ (.A(net766),
    .B(_1439_),
    .C(_1440_),
    .Y(_1456_));
 sg13g2_nor3_1 _2367_ (.A(net680),
    .B(_1446_),
    .C(_1447_),
    .Y(_1457_));
 sg13g2_nor3_1 _2368_ (.A(net761),
    .B(_1437_),
    .C(_1438_),
    .Y(_1458_));
 sg13g2_nor3_1 _2369_ (.A(net677),
    .B(_1457_),
    .C(_1458_),
    .Y(_1459_));
 sg13g2_nor3_1 _2370_ (.A(net672),
    .B(_1456_),
    .C(_1459_),
    .Y(_1460_));
 sg13g2_nor3_1 _2371_ (.A(net772),
    .B(_1444_),
    .C(_1445_),
    .Y(_1461_));
 sg13g2_nor3_1 _2372_ (.A(net668),
    .B(_1460_),
    .C(_1461_),
    .Y(_1462_));
 sg13g2_nand3_1 _2373_ (.B(_1380_),
    .C(_1381_),
    .A(net765),
    .Y(_1463_));
 sg13g2_nand3_1 _2374_ (.B(_1448_),
    .C(_1449_),
    .A(net676),
    .Y(_1464_));
 sg13g2_nand3_1 _2375_ (.B(_1448_),
    .C(_1449_),
    .A(net765),
    .Y(_1465_));
 sg13g2_o21ai_1 _2376_ (.B1(net677),
    .Y(_1466_),
    .A1(_1457_),
    .A2(_1458_));
 sg13g2_nand3_1 _2377_ (.B(_1465_),
    .C(_1466_),
    .A(net671),
    .Y(_1467_));
 sg13g2_nand3_1 _2378_ (.B(_1463_),
    .C(_1464_),
    .A(net770),
    .Y(_1468_));
 sg13g2_a21oi_1 _2379_ (.A1(net764),
    .A2(_1450_),
    .Y(_1469_),
    .B1(net772));
 sg13g2_a21oi_1 _2380_ (.A1(_1451_),
    .A2(_1452_),
    .Y(_1470_),
    .B1(net672));
 sg13g2_nor3_1 _2381_ (.A(net778),
    .B(_1469_),
    .C(_1470_),
    .Y(_1471_));
 sg13g2_nor3_1 _2382_ (.A(net668),
    .B(_1453_),
    .C(_1454_),
    .Y(_1472_));
 sg13g2_nor3_1 _2383_ (.A(net663),
    .B(_1455_),
    .C(_1462_),
    .Y(_1473_));
 sg13g2_nor3_1 _2384_ (.A(net784),
    .B(_1471_),
    .C(_1472_),
    .Y(_1474_));
 sg13g2_o21ai_1 _2385_ (.B1(net663),
    .Y(_1475_),
    .A1(_1455_),
    .A2(_1462_));
 sg13g2_o21ai_1 _2386_ (.B1(net672),
    .Y(_1476_),
    .A1(_1456_),
    .A2(_1459_));
 sg13g2_nand3_1 _2387_ (.B(_1465_),
    .C(_1466_),
    .A(net770),
    .Y(_1477_));
 sg13g2_nand3_1 _2388_ (.B(_1476_),
    .C(_1477_),
    .A(net776),
    .Y(_1478_));
 sg13g2_o21ai_1 _2389_ (.B1(net668),
    .Y(_1479_),
    .A1(_1460_),
    .A2(_1461_));
 sg13g2_nand3_1 _2390_ (.B(_1478_),
    .C(_1479_),
    .A(net782),
    .Y(_1480_));
 sg13g2_nand3_1 _2391_ (.B(_1475_),
    .C(_1480_),
    .A(net790),
    .Y(_1481_));
 sg13g2_o21ai_1 _2392_ (.B1(net658),
    .Y(_1482_),
    .A1(_1473_),
    .A2(_1474_));
 sg13g2_nand3_1 _2393_ (.B(_1463_),
    .C(_1464_),
    .A(net670),
    .Y(_1483_));
 sg13g2_nand3_1 _2394_ (.B(_1382_),
    .C(_1383_),
    .A(net770),
    .Y(_1484_));
 sg13g2_nand3_1 _2395_ (.B(_1483_),
    .C(_1484_),
    .A(net776),
    .Y(_1485_));
 sg13g2_nand3_1 _2396_ (.B(_1467_),
    .C(_1468_),
    .A(net666),
    .Y(_1486_));
 sg13g2_nand3_1 _2397_ (.B(_1467_),
    .C(_1468_),
    .A(net776),
    .Y(_1487_));
 sg13g2_nand3_1 _2398_ (.B(_1476_),
    .C(_1477_),
    .A(net666),
    .Y(_1488_));
 sg13g2_nand3_1 _2399_ (.B(_1487_),
    .C(_1488_),
    .A(net661),
    .Y(_1489_));
 sg13g2_nand3_1 _2400_ (.B(_1485_),
    .C(_1486_),
    .A(net783),
    .Y(_1490_));
 sg13g2_nand3_1 _2401_ (.B(_1489_),
    .C(_1490_),
    .A(net790),
    .Y(_1491_));
 sg13g2_nand3_1 _2402_ (.B(_1478_),
    .C(_1479_),
    .A(net661),
    .Y(_1492_));
 sg13g2_nand3_1 _2403_ (.B(_1487_),
    .C(_1488_),
    .A(net782),
    .Y(_1493_));
 sg13g2_nand3_1 _2404_ (.B(_1492_),
    .C(_1493_),
    .A(net656),
    .Y(_1494_));
 sg13g2_a21oi_1 _2405_ (.A1(_1481_),
    .A2(_1482_),
    .Y(_1495_),
    .B1(net649));
 sg13g2_o21ai_1 _2406_ (.B1(net789),
    .Y(_1496_),
    .A1(_1473_),
    .A2(_1474_));
 sg13g2_nand3_1 _2407_ (.B(net772),
    .C(_1450_),
    .A(net764),
    .Y(_1497_));
 sg13g2_nand2_1 _2408_ (.Y(_1498_),
    .A(net668),
    .B(_1497_));
 sg13g2_o21ai_1 _2409_ (.B1(net778),
    .Y(_1499_),
    .A1(_1469_),
    .A2(_1470_));
 sg13g2_nand3_1 _2410_ (.B(_1498_),
    .C(_1499_),
    .A(net663),
    .Y(_1500_));
 sg13g2_o21ai_1 _2411_ (.B1(net784),
    .Y(_1501_),
    .A1(_1471_),
    .A2(_1472_));
 sg13g2_nand3_1 _2412_ (.B(_1500_),
    .C(_1501_),
    .A(net658),
    .Y(_1502_));
 sg13g2_a21oi_1 _2413_ (.A1(_1496_),
    .A2(_1502_),
    .Y(_1503_),
    .B1(net798));
 sg13g2_nand3_1 _2414_ (.B(_1384_),
    .C(_1385_),
    .A(net776),
    .Y(_1504_));
 sg13g2_nand3_1 _2415_ (.B(_1483_),
    .C(_1484_),
    .A(net666),
    .Y(_1505_));
 sg13g2_nand3_1 _2416_ (.B(_1485_),
    .C(_1486_),
    .A(net661),
    .Y(_1506_));
 sg13g2_nand3_1 _2417_ (.B(_1504_),
    .C(_1505_),
    .A(net782),
    .Y(_1507_));
 sg13g2_nand3_1 _2418_ (.B(_1506_),
    .C(_1507_),
    .A(net790),
    .Y(_1508_));
 sg13g2_nand3_1 _2419_ (.B(_1489_),
    .C(_1490_),
    .A(net656),
    .Y(_1509_));
 sg13g2_nand3_1 _2420_ (.B(_1491_),
    .C(_1494_),
    .A(net651),
    .Y(_1510_));
 sg13g2_nand3_1 _2421_ (.B(_1508_),
    .C(_1509_),
    .A(net796),
    .Y(_1511_));
 sg13g2_nand3_1 _2422_ (.B(_1510_),
    .C(_1511_),
    .A(net804),
    .Y(_1512_));
 sg13g2_nand3_1 _2423_ (.B(_1492_),
    .C(_1493_),
    .A(net790),
    .Y(_1513_));
 sg13g2_nand3_1 _2424_ (.B(_1475_),
    .C(_1480_),
    .A(net656),
    .Y(_1514_));
 sg13g2_nand3_1 _2425_ (.B(_1513_),
    .C(_1514_),
    .A(net652),
    .Y(_1515_));
 sg13g2_nand3_1 _2426_ (.B(_1491_),
    .C(_1494_),
    .A(net796),
    .Y(_1516_));
 sg13g2_nand3_1 _2427_ (.B(_1515_),
    .C(_1516_),
    .A(net643),
    .Y(_1517_));
 sg13g2_nand3_1 _2428_ (.B(_1515_),
    .C(_1516_),
    .A(net804),
    .Y(_1518_));
 sg13g2_nand3_1 _2429_ (.B(_1481_),
    .C(_1482_),
    .A(net652),
    .Y(_1519_));
 sg13g2_nand3_1 _2430_ (.B(_1513_),
    .C(_1514_),
    .A(net796),
    .Y(_1520_));
 sg13g2_nand3_1 _2431_ (.B(_1519_),
    .C(_1520_),
    .A(net643),
    .Y(_1521_));
 sg13g2_nand3_1 _2432_ (.B(_1518_),
    .C(_1521_),
    .A(net637),
    .Y(_1522_));
 sg13g2_nand3_1 _2433_ (.B(_1512_),
    .C(_1517_),
    .A(net810),
    .Y(_1523_));
 sg13g2_nand3_1 _2434_ (.B(_1522_),
    .C(_1523_),
    .A(net818),
    .Y(_1524_));
 sg13g2_nand3_1 _2435_ (.B(_1519_),
    .C(_1520_),
    .A(net804),
    .Y(_1525_));
 sg13g2_nor3_1 _2436_ (.A(net663),
    .B(_1471_),
    .C(_1472_),
    .Y(_1526_));
 sg13g2_a21oi_1 _2437_ (.A1(_1498_),
    .A2(_1499_),
    .Y(_1527_),
    .B1(net784));
 sg13g2_nor3_1 _2438_ (.A(net789),
    .B(_1526_),
    .C(_1527_),
    .Y(_1528_));
 sg13g2_nor3_1 _2439_ (.A(net658),
    .B(_1473_),
    .C(_1474_),
    .Y(_1529_));
 sg13g2_o21ai_1 _2440_ (.B1(net649),
    .Y(_1530_),
    .A1(_1528_),
    .A2(_1529_));
 sg13g2_nand3_1 _2441_ (.B(_1481_),
    .C(_1482_),
    .A(net798),
    .Y(_1531_));
 sg13g2_nand3_1 _2442_ (.B(_1530_),
    .C(_1531_),
    .A(net645),
    .Y(_1532_));
 sg13g2_nand2_1 _2443_ (.Y(_1533_),
    .A(_1525_),
    .B(_1532_));
 sg13g2_nand3_1 _2444_ (.B(_1525_),
    .C(_1532_),
    .A(net637),
    .Y(_1534_));
 sg13g2_nand3_1 _2445_ (.B(_1518_),
    .C(_1521_),
    .A(net810),
    .Y(_1535_));
 sg13g2_nand3_1 _2446_ (.B(_1534_),
    .C(_1535_),
    .A(net630),
    .Y(_1536_));
 sg13g2_and2_1 _2447_ (.A(_1524_),
    .B(_1536_),
    .X(_1537_));
 sg13g2_nand3_1 _2448_ (.B(_1500_),
    .C(_1501_),
    .A(net792),
    .Y(_1538_));
 sg13g2_nor2_1 _2449_ (.A(net668),
    .B(_1497_),
    .Y(_1539_));
 sg13g2_nor2_1 _2450_ (.A(net784),
    .B(_1539_),
    .Y(_1540_));
 sg13g2_a21oi_1 _2451_ (.A1(_1498_),
    .A2(_1499_),
    .Y(_1541_),
    .B1(net663));
 sg13g2_o21ai_1 _2452_ (.B1(net658),
    .Y(_1542_),
    .A1(_1540_),
    .A2(_1541_));
 sg13g2_nand3_1 _2453_ (.B(_1538_),
    .C(_1542_),
    .A(net650),
    .Y(_1543_));
 sg13g2_nand3_1 _2454_ (.B(_1496_),
    .C(_1502_),
    .A(net798),
    .Y(_1544_));
 sg13g2_a21oi_1 _2455_ (.A1(_1543_),
    .A2(_1544_),
    .Y(_1545_),
    .B1(net803));
 sg13g2_nor3_1 _2456_ (.A(net645),
    .B(_1495_),
    .C(_1503_),
    .Y(_1546_));
 sg13g2_and3_1 _2457_ (.X(_1547_),
    .A(net818),
    .B(_1534_),
    .C(_1535_));
 sg13g2_nand3_1 _2458_ (.B(_1530_),
    .C(_1531_),
    .A(net803),
    .Y(_1548_));
 sg13g2_nor3_1 _2459_ (.A(net650),
    .B(_1528_),
    .C(_1529_),
    .Y(_1549_));
 sg13g2_nor3_1 _2460_ (.A(net789),
    .B(_1540_),
    .C(_1541_),
    .Y(_1550_));
 sg13g2_nor3_1 _2461_ (.A(net658),
    .B(_1526_),
    .C(_1527_),
    .Y(_1551_));
 sg13g2_nor3_1 _2462_ (.A(net798),
    .B(_1550_),
    .C(_1551_),
    .Y(_1552_));
 sg13g2_nor2_1 _2463_ (.A(_1549_),
    .B(_1552_),
    .Y(_1553_));
 sg13g2_o21ai_1 _2464_ (.B1(_1548_),
    .Y(_1554_),
    .A1(net803),
    .A2(_1553_));
 sg13g2_mux2_1 _2465_ (.A0(_1533_),
    .A1(_1554_),
    .S(net636),
    .X(_1555_));
 sg13g2_a21oi_1 _2466_ (.A1(net630),
    .A2(_1555_),
    .Y(_1556_),
    .B1(_1547_));
 sg13g2_a21oi_1 _2467_ (.A1(\ayayayayayaya.b[28] ),
    .A2(net623),
    .Y(_1557_),
    .B1(_0611_));
 sg13g2_a22oi_1 _2468_ (.Y(_1558_),
    .B1(net615),
    .B2(net718),
    .A2(net620),
    .A1(net749));
 sg13g2_nand2_1 _2469_ (.Y(_1559_),
    .A(net842),
    .B(\a[24] ));
 sg13g2_o21ai_1 _2470_ (.B1(\a[25] ),
    .Y(_1560_),
    .A1(net838),
    .A2(_1559_));
 sg13g2_a21oi_1 _2471_ (.A1(net834),
    .A2(_1559_),
    .Y(_1561_),
    .B1(_1560_));
 sg13g2_o21ai_1 _2472_ (.B1(net607),
    .Y(_1562_),
    .A1(\a[25] ),
    .A2(net834));
 sg13g2_a21oi_1 _2473_ (.A1(\a[24] ),
    .A2(_1562_),
    .Y(_1563_),
    .B1(_1561_));
 sg13g2_nand3_1 _2474_ (.B(_1558_),
    .C(_1563_),
    .A(_1557_),
    .Y(_1564_));
 sg13g2_a21oi_1 _2475_ (.A1(_1003_),
    .A2(_1004_),
    .Y(_1565_),
    .B1(net602));
 sg13g2_or2_1 _2476_ (.X(_1566_),
    .B(_1565_),
    .A(_1564_));
 sg13g2_a221oi_1 _2477_ (.B2(net595),
    .C1(_1566_),
    .B1(_1556_),
    .A1(net601),
    .Y(_1567_),
    .A2(_1537_));
 sg13g2_nand3b_1 _2478_ (.B(net843),
    .C(_1427_),
    .Y(_1568_),
    .A_N(_1567_));
 sg13g2_a21oi_1 _2479_ (.A1(_1339_),
    .A2(_1340_),
    .Y(_1569_),
    .B1(net745));
 sg13g2_or3_1 _2480_ (.A(net741),
    .B(_1337_),
    .C(_1338_),
    .X(_1570_));
 sg13g2_nand2_1 _2481_ (.Y(_1571_),
    .A(net824),
    .B(net741));
 sg13g2_and3_1 _2482_ (.X(_1572_),
    .A(net745),
    .B(_1570_),
    .C(_1571_));
 sg13g2_o21ai_1 _2483_ (.B1(net748),
    .Y(_1573_),
    .A1(_1569_),
    .A2(_1572_));
 sg13g2_nand3_1 _2484_ (.B(_1341_),
    .C(_1342_),
    .A(net692),
    .Y(_1574_));
 sg13g2_nand3_1 _2485_ (.B(_1343_),
    .C(_1344_),
    .A(net688),
    .Y(_1575_));
 sg13g2_nand3_1 _2486_ (.B(_1573_),
    .C(_1574_),
    .A(net749),
    .Y(_1576_));
 sg13g2_nor2_1 _2487_ (.A(\a[14] ),
    .B(net696),
    .Y(_1577_));
 sg13g2_a21oi_1 _2488_ (.A1(net696),
    .A2(_1571_),
    .Y(_1578_),
    .B1(_1577_));
 sg13g2_nor2_1 _2489_ (.A(net692),
    .B(_1578_),
    .Y(_1579_));
 sg13g2_o21ai_1 _2490_ (.B1(_1579_),
    .Y(_1580_),
    .A1(_1570_),
    .A2(_1577_));
 sg13g2_o21ai_1 _2491_ (.B1(net692),
    .Y(_1581_),
    .A1(_1569_),
    .A2(_1572_));
 sg13g2_nand3_1 _2492_ (.B(_1573_),
    .C(_1574_),
    .A(net688),
    .Y(_1582_));
 sg13g2_nand3_1 _2493_ (.B(_1580_),
    .C(_1581_),
    .A(net749),
    .Y(_1583_));
 sg13g2_nand3_1 _2494_ (.B(_1582_),
    .C(_1583_),
    .A(net753),
    .Y(_1584_));
 sg13g2_nand3_1 _2495_ (.B(_1575_),
    .C(_1576_),
    .A(net685),
    .Y(_1585_));
 sg13g2_nand3_1 _2496_ (.B(_1575_),
    .C(_1576_),
    .A(net754),
    .Y(_1586_));
 sg13g2_nand3_1 _2497_ (.B(_1345_),
    .C(_1346_),
    .A(net685),
    .Y(_1587_));
 sg13g2_nand3_1 _2498_ (.B(_1586_),
    .C(_1587_),
    .A(net681),
    .Y(_1588_));
 sg13g2_nand3_1 _2499_ (.B(_1584_),
    .C(_1585_),
    .A(net759),
    .Y(_1589_));
 sg13g2_a21oi_1 _2500_ (.A1(_1580_),
    .A2(_1581_),
    .Y(_1590_),
    .B1(net749));
 sg13g2_nor2_1 _2501_ (.A(\a[13] ),
    .B(net692),
    .Y(_1591_));
 sg13g2_nor3_1 _2502_ (.A(_1570_),
    .B(_1577_),
    .C(_1591_),
    .Y(_1592_));
 sg13g2_nor2_1 _2503_ (.A(net748),
    .B(_1578_),
    .Y(_1593_));
 sg13g2_nor2_1 _2504_ (.A(_1591_),
    .B(_1593_),
    .Y(_1594_));
 sg13g2_nor3_1 _2505_ (.A(net688),
    .B(_1592_),
    .C(_1594_),
    .Y(_1595_));
 sg13g2_o21ai_1 _2506_ (.B1(net753),
    .Y(_1596_),
    .A1(_1590_),
    .A2(_1595_));
 sg13g2_nand3_1 _2507_ (.B(_1582_),
    .C(_1583_),
    .A(net685),
    .Y(_1597_));
 sg13g2_nand3_1 _2508_ (.B(_1584_),
    .C(_1585_),
    .A(net681),
    .Y(_1598_));
 sg13g2_nand3_1 _2509_ (.B(_1596_),
    .C(_1597_),
    .A(net759),
    .Y(_1599_));
 sg13g2_nand3_1 _2510_ (.B(_1598_),
    .C(_1599_),
    .A(net763),
    .Y(_1600_));
 sg13g2_nand3_1 _2511_ (.B(_1588_),
    .C(_1589_),
    .A(net675),
    .Y(_1601_));
 sg13g2_nand3_1 _2512_ (.B(_1347_),
    .C(_1348_),
    .A(net681),
    .Y(_1602_));
 sg13g2_nand3_1 _2513_ (.B(_1586_),
    .C(_1587_),
    .A(net759),
    .Y(_1603_));
 sg13g2_nand3_1 _2514_ (.B(_1588_),
    .C(_1589_),
    .A(net764),
    .Y(_1604_));
 sg13g2_nand3_1 _2515_ (.B(_1602_),
    .C(_1603_),
    .A(net675),
    .Y(_1605_));
 sg13g2_nand3_1 _2516_ (.B(_1604_),
    .C(_1605_),
    .A(net673),
    .Y(_1606_));
 sg13g2_nand3_1 _2517_ (.B(_1600_),
    .C(_1601_),
    .A(net769),
    .Y(_1607_));
 sg13g2_nor2_1 _2518_ (.A(\a[12] ),
    .B(net688),
    .Y(_1608_));
 sg13g2_nand2b_1 _2519_ (.Y(_1609_),
    .B(_1592_),
    .A_N(_1608_));
 sg13g2_nor2_1 _2520_ (.A(net749),
    .B(_1594_),
    .Y(_1610_));
 sg13g2_nor2_1 _2521_ (.A(_1608_),
    .B(_1610_),
    .Y(_1611_));
 sg13g2_nor2_1 _2522_ (.A(net685),
    .B(_1611_),
    .Y(_1612_));
 sg13g2_nand2_1 _2523_ (.Y(_1613_),
    .A(_1609_),
    .B(_1612_));
 sg13g2_o21ai_1 _2524_ (.B1(net685),
    .Y(_1614_),
    .A1(_1590_),
    .A2(_1595_));
 sg13g2_nand3_1 _2525_ (.B(_1596_),
    .C(_1597_),
    .A(net681),
    .Y(_1615_));
 sg13g2_nand3_1 _2526_ (.B(_1613_),
    .C(_1614_),
    .A(net758),
    .Y(_1616_));
 sg13g2_nand3_1 _2527_ (.B(_1615_),
    .C(_1616_),
    .A(net763),
    .Y(_1617_));
 sg13g2_nand3_1 _2528_ (.B(_1598_),
    .C(_1599_),
    .A(net675),
    .Y(_1618_));
 sg13g2_nand3_1 _2529_ (.B(_1600_),
    .C(_1601_),
    .A(net669),
    .Y(_1619_));
 sg13g2_nand3_1 _2530_ (.B(_1617_),
    .C(_1618_),
    .A(net769),
    .Y(_1620_));
 sg13g2_nand3_1 _2531_ (.B(_1619_),
    .C(_1620_),
    .A(net775),
    .Y(_1621_));
 sg13g2_nand3_1 _2532_ (.B(_1606_),
    .C(_1607_),
    .A(net665),
    .Y(_1622_));
 sg13g2_nand3_1 _2533_ (.B(_1602_),
    .C(_1603_),
    .A(net764),
    .Y(_1623_));
 sg13g2_nand3_1 _2534_ (.B(_1349_),
    .C(_1350_),
    .A(net677),
    .Y(_1624_));
 sg13g2_nand3_1 _2535_ (.B(_1623_),
    .C(_1624_),
    .A(net672),
    .Y(_1625_));
 sg13g2_nand3_1 _2536_ (.B(_1604_),
    .C(_1605_),
    .A(net769),
    .Y(_1626_));
 sg13g2_nand3_1 _2537_ (.B(_1606_),
    .C(_1607_),
    .A(net775),
    .Y(_1627_));
 sg13g2_nand3_1 _2538_ (.B(_1625_),
    .C(_1626_),
    .A(net668),
    .Y(_1628_));
 sg13g2_nand3_1 _2539_ (.B(_1627_),
    .C(_1628_),
    .A(net660),
    .Y(_1629_));
 sg13g2_nand3_1 _2540_ (.B(_1621_),
    .C(_1622_),
    .A(net781),
    .Y(_1630_));
 sg13g2_a21oi_1 _2541_ (.A1(_1613_),
    .A2(_1614_),
    .Y(_1631_),
    .B1(net758));
 sg13g2_nand2b_2 _2542_ (.Y(_1632_),
    .B(net754),
    .A_N(\a[11] ));
 sg13g2_nand2b_1 _2543_ (.Y(_1633_),
    .B(_1632_),
    .A_N(_1609_));
 sg13g2_o21ai_1 _2544_ (.B1(_1632_),
    .Y(_1634_),
    .A1(net753),
    .A2(_1611_));
 sg13g2_and3_1 _2545_ (.X(_1635_),
    .A(net758),
    .B(_1633_),
    .C(_1634_));
 sg13g2_o21ai_1 _2546_ (.B1(net763),
    .Y(_1636_),
    .A1(_1631_),
    .A2(_1635_));
 sg13g2_nand3_1 _2547_ (.B(_1615_),
    .C(_1616_),
    .A(net674),
    .Y(_1637_));
 sg13g2_nand3_1 _2548_ (.B(_1617_),
    .C(_1618_),
    .A(net673),
    .Y(_1638_));
 sg13g2_nand3_1 _2549_ (.B(_1636_),
    .C(_1637_),
    .A(net769),
    .Y(_1639_));
 sg13g2_nand3_1 _2550_ (.B(_1638_),
    .C(_1639_),
    .A(net775),
    .Y(_1640_));
 sg13g2_nand3_1 _2551_ (.B(_1619_),
    .C(_1620_),
    .A(net665),
    .Y(_1641_));
 sg13g2_nand3_1 _2552_ (.B(_1621_),
    .C(_1622_),
    .A(net660),
    .Y(_1642_));
 sg13g2_nand3_1 _2553_ (.B(_1640_),
    .C(_1641_),
    .A(net781),
    .Y(_1643_));
 sg13g2_nand3_1 _2554_ (.B(_1642_),
    .C(_1643_),
    .A(net787),
    .Y(_1644_));
 sg13g2_nand3_1 _2555_ (.B(_1629_),
    .C(_1630_),
    .A(net655),
    .Y(_1645_));
 sg13g2_nand3_1 _2556_ (.B(_1351_),
    .C(_1352_),
    .A(net672),
    .Y(_1646_));
 sg13g2_nand3_1 _2557_ (.B(_1623_),
    .C(_1624_),
    .A(net772),
    .Y(_1647_));
 sg13g2_nand3_1 _2558_ (.B(_1625_),
    .C(_1626_),
    .A(net778),
    .Y(_1648_));
 sg13g2_nand3_1 _2559_ (.B(_1646_),
    .C(_1647_),
    .A(net668),
    .Y(_1649_));
 sg13g2_nand3_1 _2560_ (.B(_1648_),
    .C(_1649_),
    .A(net663),
    .Y(_1650_));
 sg13g2_nand3_1 _2561_ (.B(_1627_),
    .C(_1628_),
    .A(net781),
    .Y(_1651_));
 sg13g2_nand3_1 _2562_ (.B(_1629_),
    .C(_1630_),
    .A(net787),
    .Y(_1652_));
 sg13g2_nand3_1 _2563_ (.B(_1650_),
    .C(_1651_),
    .A(net658),
    .Y(_1653_));
 sg13g2_nand3_1 _2564_ (.B(_1652_),
    .C(_1653_),
    .A(net649),
    .Y(_1654_));
 sg13g2_nand3_1 _2565_ (.B(_1644_),
    .C(_1645_),
    .A(net794),
    .Y(_1655_));
 sg13g2_nand2b_2 _2566_ (.Y(_1656_),
    .B(net762),
    .A_N(\a[10] ));
 sg13g2_nand2b_1 _2567_ (.Y(_1657_),
    .B(_1656_),
    .A_N(_1633_));
 sg13g2_nand2_1 _2568_ (.Y(_1658_),
    .A(net681),
    .B(_1634_));
 sg13g2_and2_1 _2569_ (.A(_1656_),
    .B(_1658_),
    .X(_1659_));
 sg13g2_nor2_1 _2570_ (.A(net674),
    .B(_1659_),
    .Y(_1660_));
 sg13g2_nand2_1 _2571_ (.Y(_1661_),
    .A(_1657_),
    .B(_1660_));
 sg13g2_o21ai_1 _2572_ (.B1(net674),
    .Y(_1662_),
    .A1(_1631_),
    .A2(_1635_));
 sg13g2_nand3_1 _2573_ (.B(_1636_),
    .C(_1637_),
    .A(net669),
    .Y(_1663_));
 sg13g2_nand3_1 _2574_ (.B(_1661_),
    .C(_1662_),
    .A(net768),
    .Y(_1664_));
 sg13g2_nand3_1 _2575_ (.B(_1663_),
    .C(_1664_),
    .A(net775),
    .Y(_1665_));
 sg13g2_nand3_1 _2576_ (.B(_1638_),
    .C(_1639_),
    .A(net665),
    .Y(_1666_));
 sg13g2_nand3_1 _2577_ (.B(_1640_),
    .C(_1641_),
    .A(net660),
    .Y(_1667_));
 sg13g2_nand3_1 _2578_ (.B(_1665_),
    .C(_1666_),
    .A(net781),
    .Y(_1668_));
 sg13g2_nand3_1 _2579_ (.B(_1667_),
    .C(_1668_),
    .A(net787),
    .Y(_1669_));
 sg13g2_nand3_1 _2580_ (.B(_1642_),
    .C(_1643_),
    .A(net655),
    .Y(_1670_));
 sg13g2_nand3_1 _2581_ (.B(_1644_),
    .C(_1645_),
    .A(net648),
    .Y(_1671_));
 sg13g2_nand3_1 _2582_ (.B(_1669_),
    .C(_1670_),
    .A(net794),
    .Y(_1672_));
 sg13g2_nand3_1 _2583_ (.B(_1671_),
    .C(_1672_),
    .A(net800),
    .Y(_1673_));
 sg13g2_nand3_1 _2584_ (.B(_1654_),
    .C(_1655_),
    .A(net642),
    .Y(_1674_));
 sg13g2_nand3_1 _2585_ (.B(_1646_),
    .C(_1647_),
    .A(net778),
    .Y(_1675_));
 sg13g2_nand3_1 _2586_ (.B(_1353_),
    .C(_1354_),
    .A(net666),
    .Y(_1676_));
 sg13g2_nand3_1 _2587_ (.B(_1675_),
    .C(_1676_),
    .A(net663),
    .Y(_1677_));
 sg13g2_nand3_1 _2588_ (.B(_1648_),
    .C(_1649_),
    .A(net784),
    .Y(_0064_));
 sg13g2_nand3_1 _2589_ (.B(_1650_),
    .C(_1651_),
    .A(net789),
    .Y(_0065_));
 sg13g2_nand3_1 _2590_ (.B(_1677_),
    .C(_0064_),
    .A(net658),
    .Y(_0066_));
 sg13g2_nand3_1 _2591_ (.B(_0065_),
    .C(_0066_),
    .A(net649),
    .Y(_0067_));
 sg13g2_nand3_1 _2592_ (.B(_1652_),
    .C(_1653_),
    .A(net798),
    .Y(_0068_));
 sg13g2_nand3_1 _2593_ (.B(_1654_),
    .C(_1655_),
    .A(net801),
    .Y(_0069_));
 sg13g2_nand3_1 _2594_ (.B(_0067_),
    .C(_0068_),
    .A(net645),
    .Y(_0070_));
 sg13g2_nand3_1 _2595_ (.B(_0069_),
    .C(_0070_),
    .A(net636),
    .Y(_0071_));
 sg13g2_nand3_1 _2596_ (.B(_1673_),
    .C(_1674_),
    .A(net807),
    .Y(_0072_));
 sg13g2_a21oi_1 _2597_ (.A1(_1661_),
    .A2(_1662_),
    .Y(_0073_),
    .B1(net768));
 sg13g2_a21oi_1 _2598_ (.A1(_0654_),
    .A2(net763),
    .Y(_0074_),
    .B1(_1657_));
 sg13g2_nor2_1 _2599_ (.A(net763),
    .B(_1659_),
    .Y(_0075_));
 sg13g2_a21oi_1 _2600_ (.A1(_0654_),
    .A2(net763),
    .Y(_0076_),
    .B1(_0075_));
 sg13g2_nor3_1 _2601_ (.A(net669),
    .B(_0074_),
    .C(_0076_),
    .Y(_0077_));
 sg13g2_o21ai_1 _2602_ (.B1(net774),
    .Y(_0078_),
    .A1(_0073_),
    .A2(_0077_));
 sg13g2_nand3_1 _2603_ (.B(_1663_),
    .C(_1664_),
    .A(net664),
    .Y(_0079_));
 sg13g2_nand3_1 _2604_ (.B(_1665_),
    .C(_1666_),
    .A(net660),
    .Y(_0080_));
 sg13g2_nand3_1 _2605_ (.B(_0078_),
    .C(_0079_),
    .A(net780),
    .Y(_0081_));
 sg13g2_nand3_1 _2606_ (.B(_0080_),
    .C(_0081_),
    .A(net787),
    .Y(_0082_));
 sg13g2_nand3_1 _2607_ (.B(_1667_),
    .C(_1668_),
    .A(net655),
    .Y(_0083_));
 sg13g2_nand3_1 _2608_ (.B(_1669_),
    .C(_1670_),
    .A(net648),
    .Y(_0084_));
 sg13g2_nand3_1 _2609_ (.B(_0082_),
    .C(_0083_),
    .A(net794),
    .Y(_0085_));
 sg13g2_nand3_1 _2610_ (.B(_0084_),
    .C(_0085_),
    .A(net801),
    .Y(_0086_));
 sg13g2_nand3_1 _2611_ (.B(_1671_),
    .C(_1672_),
    .A(net642),
    .Y(_0087_));
 sg13g2_nand3_1 _2612_ (.B(_1673_),
    .C(_1674_),
    .A(net635),
    .Y(_0088_));
 sg13g2_nand3_1 _2613_ (.B(_0086_),
    .C(_0087_),
    .A(net807),
    .Y(_0089_));
 sg13g2_nand3_1 _2614_ (.B(_0088_),
    .C(_0089_),
    .A(net814),
    .Y(_0090_));
 sg13g2_nand3_1 _2615_ (.B(_0071_),
    .C(_0072_),
    .A(net629),
    .Y(_0091_));
 sg13g2_nand3_1 _2616_ (.B(_0090_),
    .C(_0091_),
    .A(net594),
    .Y(_0092_));
 sg13g2_nand2b_1 _2617_ (.Y(_0093_),
    .B(net769),
    .A_N(net825));
 sg13g2_and2_1 _2618_ (.A(_0074_),
    .B(_0093_),
    .X(_0094_));
 sg13g2_mux2_1 _2619_ (.A0(net825),
    .A1(_0076_),
    .S(net669),
    .X(_0095_));
 sg13g2_nor2_1 _2620_ (.A(net665),
    .B(_0095_),
    .Y(_0096_));
 sg13g2_nand2b_1 _2621_ (.Y(_0097_),
    .B(_0096_),
    .A_N(_0094_));
 sg13g2_o21ai_1 _2622_ (.B1(net664),
    .Y(_0098_),
    .A1(_0073_),
    .A2(_0077_));
 sg13g2_nand3_1 _2623_ (.B(_0078_),
    .C(_0079_),
    .A(net659),
    .Y(_0099_));
 sg13g2_nand3_1 _2624_ (.B(_0097_),
    .C(_0098_),
    .A(net781),
    .Y(_0100_));
 sg13g2_nand3_1 _2625_ (.B(_0099_),
    .C(_0100_),
    .A(net786),
    .Y(_0101_));
 sg13g2_nand3_1 _2626_ (.B(_0080_),
    .C(_0081_),
    .A(net655),
    .Y(_0102_));
 sg13g2_nand3_1 _2627_ (.B(_0082_),
    .C(_0083_),
    .A(net648),
    .Y(_0103_));
 sg13g2_nand3_1 _2628_ (.B(_0101_),
    .C(_0102_),
    .A(net793),
    .Y(_0104_));
 sg13g2_nand3_1 _2629_ (.B(_0103_),
    .C(_0104_),
    .A(net801),
    .Y(_0105_));
 sg13g2_nand3_1 _2630_ (.B(_0084_),
    .C(_0085_),
    .A(net642),
    .Y(_0106_));
 sg13g2_nand3_1 _2631_ (.B(_0086_),
    .C(_0087_),
    .A(net635),
    .Y(_0107_));
 sg13g2_nand3_1 _2632_ (.B(_0105_),
    .C(_0106_),
    .A(net807),
    .Y(_0108_));
 sg13g2_nand3_1 _2633_ (.B(_0107_),
    .C(_0108_),
    .A(net815),
    .Y(_0109_));
 sg13g2_nand3_1 _2634_ (.B(_0088_),
    .C(_0089_),
    .A(net629),
    .Y(_0110_));
 sg13g2_nand3_1 _2635_ (.B(_0109_),
    .C(_0110_),
    .A(net598),
    .Y(_0111_));
 sg13g2_and2_1 _2636_ (.A(net823),
    .B(_1423_),
    .X(_0112_));
 sg13g2_nand3_1 _2637_ (.B(net741),
    .C(net745),
    .A(net824),
    .Y(_0113_));
 sg13g2_a21oi_1 _2638_ (.A1(net692),
    .A2(_0113_),
    .Y(_0114_),
    .B1(_1579_));
 sg13g2_mux2_1 _2639_ (.A0(_1594_),
    .A1(_0114_),
    .S(net688),
    .X(_0115_));
 sg13g2_nor2_1 _2640_ (.A(net685),
    .B(_0115_),
    .Y(_0116_));
 sg13g2_nor3_1 _2641_ (.A(net692),
    .B(net749),
    .C(_0113_),
    .Y(_0117_));
 sg13g2_a21oi_1 _2642_ (.A1(net749),
    .A2(_0114_),
    .Y(_0118_),
    .B1(_0117_));
 sg13g2_a21oi_1 _2643_ (.A1(net685),
    .A2(_0118_),
    .Y(_0119_),
    .B1(_0116_));
 sg13g2_nor2_1 _2644_ (.A(net753),
    .B(_0115_),
    .Y(_0120_));
 sg13g2_nor2_1 _2645_ (.A(_1612_),
    .B(_0120_),
    .Y(_0121_));
 sg13g2_mux2_1 _2646_ (.A0(_0119_),
    .A1(_0121_),
    .S(net757),
    .X(_0122_));
 sg13g2_nand2_1 _2647_ (.Y(_0123_),
    .A(net753),
    .B(_0118_));
 sg13g2_nor3_2 _2648_ (.A(net692),
    .B(net688),
    .C(_0113_),
    .Y(_0124_));
 sg13g2_o21ai_1 _2649_ (.B1(_0123_),
    .Y(_0125_),
    .A1(net753),
    .A2(_0124_));
 sg13g2_nand2_1 _2650_ (.Y(_0126_),
    .A(net757),
    .B(_0119_));
 sg13g2_o21ai_1 _2651_ (.B1(_0126_),
    .Y(_0127_),
    .A1(net757),
    .A2(_0125_));
 sg13g2_mux2_1 _2652_ (.A0(_0122_),
    .A1(_0127_),
    .S(net674),
    .X(_0128_));
 sg13g2_nor2_1 _2653_ (.A(net757),
    .B(_0121_),
    .Y(_0129_));
 sg13g2_a21oi_1 _2654_ (.A1(net757),
    .A2(_1634_),
    .Y(_0130_),
    .B1(_0129_));
 sg13g2_mux2_1 _2655_ (.A0(_0122_),
    .A1(_0130_),
    .S(net763),
    .X(_0131_));
 sg13g2_mux2_1 _2656_ (.A0(_0128_),
    .A1(_0131_),
    .S(net768),
    .X(_0132_));
 sg13g2_a21oi_1 _2657_ (.A1(net753),
    .A2(_0124_),
    .Y(_0133_),
    .B1(net757));
 sg13g2_a21oi_1 _2658_ (.A1(net757),
    .A2(_0125_),
    .Y(_0134_),
    .B1(_0133_));
 sg13g2_mux2_1 _2659_ (.A0(_0127_),
    .A1(_0134_),
    .S(net674),
    .X(_0135_));
 sg13g2_mux2_1 _2660_ (.A0(_0128_),
    .A1(_0135_),
    .S(net669),
    .X(_0136_));
 sg13g2_mux2_1 _2661_ (.A0(_0132_),
    .A1(_0136_),
    .S(net664),
    .X(_0137_));
 sg13g2_nor2_1 _2662_ (.A(net763),
    .B(_0130_),
    .Y(_0138_));
 sg13g2_nor2_1 _2663_ (.A(_1660_),
    .B(_0138_),
    .Y(_0139_));
 sg13g2_mux2_1 _2664_ (.A0(_0131_),
    .A1(_0139_),
    .S(net768),
    .X(_0140_));
 sg13g2_mux2_1 _2665_ (.A0(_0132_),
    .A1(_0140_),
    .S(net774),
    .X(_0141_));
 sg13g2_mux2_1 _2666_ (.A0(_0137_),
    .A1(_0141_),
    .S(net780),
    .X(_0142_));
 sg13g2_nand3_1 _2667_ (.B(net757),
    .C(_0124_),
    .A(net753),
    .Y(_0143_));
 sg13g2_nand2_1 _2668_ (.Y(_0144_),
    .A(net674),
    .B(_0143_));
 sg13g2_o21ai_1 _2669_ (.B1(_0144_),
    .Y(_0145_),
    .A1(net674),
    .A2(_0134_));
 sg13g2_nand2_1 _2670_ (.Y(_0146_),
    .A(net768),
    .B(_0135_));
 sg13g2_o21ai_1 _2671_ (.B1(_0146_),
    .Y(_0147_),
    .A1(net768),
    .A2(_0145_));
 sg13g2_mux2_1 _2672_ (.A0(_0136_),
    .A1(_0147_),
    .S(net664),
    .X(_0148_));
 sg13g2_mux2_1 _2673_ (.A0(_0137_),
    .A1(_0148_),
    .S(net659),
    .X(_0149_));
 sg13g2_mux2_1 _2674_ (.A0(_0142_),
    .A1(_0149_),
    .S(net654),
    .X(_0150_));
 sg13g2_mux2_1 _2675_ (.A0(_0076_),
    .A1(_0139_),
    .S(net669),
    .X(_0151_));
 sg13g2_mux2_1 _2676_ (.A0(_0140_),
    .A1(_0151_),
    .S(net774),
    .X(_0152_));
 sg13g2_mux2_1 _2677_ (.A0(_0141_),
    .A1(_0152_),
    .S(net780),
    .X(_0153_));
 sg13g2_mux2_1 _2678_ (.A0(_0142_),
    .A1(_0153_),
    .S(net786),
    .X(_0154_));
 sg13g2_mux2_1 _2679_ (.A0(_0150_),
    .A1(_0154_),
    .S(net793),
    .X(_0155_));
 sg13g2_nor2_1 _2680_ (.A(net664),
    .B(_0147_),
    .Y(_0156_));
 sg13g2_nor2_1 _2681_ (.A(net674),
    .B(_0143_),
    .Y(_0157_));
 sg13g2_nor2_1 _2682_ (.A(net669),
    .B(_0145_),
    .Y(_0158_));
 sg13g2_a21oi_1 _2683_ (.A1(net669),
    .A2(_0157_),
    .Y(_0159_),
    .B1(_0158_));
 sg13g2_a21oi_1 _2684_ (.A1(net664),
    .A2(_0159_),
    .Y(_0160_),
    .B1(_0156_));
 sg13g2_mux2_1 _2685_ (.A0(_0148_),
    .A1(_0160_),
    .S(net659),
    .X(_0161_));
 sg13g2_mux2_1 _2686_ (.A0(_0149_),
    .A1(_0161_),
    .S(net654),
    .X(_0162_));
 sg13g2_mux2_1 _2687_ (.A0(_0150_),
    .A1(_0162_),
    .S(net646),
    .X(_0163_));
 sg13g2_mux2_1 _2688_ (.A0(_0155_),
    .A1(_0163_),
    .S(net640),
    .X(_0164_));
 sg13g2_nor2_1 _2689_ (.A(net774),
    .B(_0151_),
    .Y(_0165_));
 sg13g2_nor2_1 _2690_ (.A(_0096_),
    .B(_0165_),
    .Y(_0166_));
 sg13g2_mux2_1 _2691_ (.A0(_0152_),
    .A1(_0166_),
    .S(net780),
    .X(_0167_));
 sg13g2_mux2_1 _2692_ (.A0(_0153_),
    .A1(_0167_),
    .S(net786),
    .X(_0168_));
 sg13g2_mux2_1 _2693_ (.A0(_0154_),
    .A1(_0168_),
    .S(net793),
    .X(_0169_));
 sg13g2_mux2_1 _2694_ (.A0(_0155_),
    .A1(_0169_),
    .S(net800),
    .X(_0170_));
 sg13g2_mux2_1 _2695_ (.A0(_0164_),
    .A1(_0170_),
    .S(net807),
    .X(_0171_));
 sg13g2_a21oi_1 _2696_ (.A1(net768),
    .A2(_0157_),
    .Y(_0172_),
    .B1(net774));
 sg13g2_a21oi_1 _2697_ (.A1(net774),
    .A2(_0159_),
    .Y(_0173_),
    .B1(_0172_));
 sg13g2_mux2_1 _2698_ (.A0(_0160_),
    .A1(_0173_),
    .S(net659),
    .X(_0174_));
 sg13g2_mux2_1 _2699_ (.A0(_0161_),
    .A1(_0174_),
    .S(net654),
    .X(_0175_));
 sg13g2_mux2_1 _2700_ (.A0(_0162_),
    .A1(_0175_),
    .S(net646),
    .X(_0176_));
 sg13g2_mux2_1 _2701_ (.A0(_0163_),
    .A1(_0176_),
    .S(net640),
    .X(_0177_));
 sg13g2_mux2_1 _2702_ (.A0(_0164_),
    .A1(_0177_),
    .S(net633),
    .X(_0178_));
 sg13g2_mux2_1 _2703_ (.A0(_0171_),
    .A1(_0178_),
    .S(net627),
    .X(_0179_));
 sg13g2_a21oi_1 _2704_ (.A1(net726),
    .A2(net623),
    .Y(_0180_),
    .B1(_0611_));
 sg13g2_a22oi_1 _2705_ (.Y(_0181_),
    .B1(net612),
    .B2(net773),
    .A2(net616),
    .A1(net795));
 sg13g2_and2_1 _2706_ (.A(net825),
    .B(net604),
    .X(_0182_));
 sg13g2_a21oi_1 _2707_ (.A1(net839),
    .A2(net825),
    .Y(_0183_),
    .B1(net833));
 sg13g2_o21ai_1 _2708_ (.B1(\a[9] ),
    .Y(_0184_),
    .A1(_0182_),
    .A2(_0183_));
 sg13g2_nor2_1 _2709_ (.A(\a[9] ),
    .B(net833),
    .Y(_0185_));
 sg13g2_o21ai_1 _2710_ (.B1(net825),
    .Y(_0186_),
    .A1(net609),
    .A2(_0185_));
 sg13g2_nand4_1 _2711_ (.B(_0181_),
    .C(_0184_),
    .A(_0180_),
    .Y(_0187_),
    .D(_0186_));
 sg13g2_nor2_1 _2712_ (.A(net823),
    .B(net603),
    .Y(_0188_));
 sg13g2_nand3_1 _2713_ (.B(net774),
    .C(_0157_),
    .A(net768),
    .Y(_0189_));
 sg13g2_nand2_1 _2714_ (.Y(_0190_),
    .A(net780),
    .B(_0173_));
 sg13g2_o21ai_1 _2715_ (.B1(_0190_),
    .Y(_0191_),
    .A1(net780),
    .A2(_0189_));
 sg13g2_mux2_1 _2716_ (.A0(_0174_),
    .A1(_0191_),
    .S(net654),
    .X(_0192_));
 sg13g2_mux2_1 _2717_ (.A0(_0175_),
    .A1(_0192_),
    .S(net646),
    .X(_0193_));
 sg13g2_mux2_1 _2718_ (.A0(_0176_),
    .A1(_0193_),
    .S(net640),
    .X(_0194_));
 sg13g2_mux2_1 _2719_ (.A0(_0177_),
    .A1(_0194_),
    .S(net633),
    .X(_0195_));
 sg13g2_mux2_1 _2720_ (.A0(_0178_),
    .A1(_0195_),
    .S(net628),
    .X(_0196_));
 sg13g2_a221oi_1 _2721_ (.B2(_0196_),
    .C1(_0187_),
    .B1(net589),
    .A1(net591),
    .Y(_0197_),
    .A2(_0179_));
 sg13g2_nand3_1 _2722_ (.B(_0111_),
    .C(_0197_),
    .A(_0092_),
    .Y(_0198_));
 sg13g2_nand2b_1 _2723_ (.Y(_0199_),
    .B(net775),
    .A_N(net826));
 sg13g2_mux2_1 _2724_ (.A0(net826),
    .A1(_0095_),
    .S(net664),
    .X(_0200_));
 sg13g2_mux2_1 _2725_ (.A0(\a[6] ),
    .A1(_0200_),
    .S(net659),
    .X(_0201_));
 sg13g2_nor2_1 _2726_ (.A(net788),
    .B(_0201_),
    .Y(_0202_));
 sg13g2_a21oi_1 _2727_ (.A1(_0643_),
    .A2(net788),
    .Y(_0203_),
    .B1(_0202_));
 sg13g2_mux2_1 _2728_ (.A0(\a[4] ),
    .A1(_0203_),
    .S(net646),
    .X(_0204_));
 sg13g2_nor2_1 _2729_ (.A(net802),
    .B(_0204_),
    .Y(_0205_));
 sg13g2_a21oi_1 _2730_ (.A1(_0632_),
    .A2(net802),
    .Y(_0206_),
    .B1(_0205_));
 sg13g2_mux2_1 _2731_ (.A0(\a[2] ),
    .A1(_0206_),
    .S(net633),
    .X(_0207_));
 sg13g2_nor2_1 _2732_ (.A(net816),
    .B(_0207_),
    .Y(_0208_));
 sg13g2_a21oi_1 _2733_ (.A1(_0621_),
    .A2(net816),
    .Y(_0209_),
    .B1(_0208_));
 sg13g2_nor2_1 _2734_ (.A(net822),
    .B(_0209_),
    .Y(_0210_));
 sg13g2_and2_1 _2735_ (.A(_0094_),
    .B(_0199_),
    .X(_0211_));
 sg13g2_o21ai_1 _2736_ (.B1(_0211_),
    .Y(_0212_),
    .A1(\a[6] ),
    .A2(net660));
 sg13g2_a21oi_1 _2737_ (.A1(_0643_),
    .A2(net788),
    .Y(_0213_),
    .B1(_0212_));
 sg13g2_o21ai_1 _2738_ (.B1(_0213_),
    .Y(_0214_),
    .A1(\a[4] ),
    .A2(net647));
 sg13g2_a21oi_1 _2739_ (.A1(_0632_),
    .A2(net802),
    .Y(_0215_),
    .B1(_0214_));
 sg13g2_o21ai_1 _2740_ (.B1(_0215_),
    .Y(_0216_),
    .A1(\a[2] ),
    .A2(net633));
 sg13g2_a21oi_1 _2741_ (.A1(_0621_),
    .A2(net816),
    .Y(_0217_),
    .B1(_0216_));
 sg13g2_nor2b_1 _2742_ (.A(_0217_),
    .B_N(_0210_),
    .Y(_0218_));
 sg13g2_nor2b_1 _2743_ (.A(net827),
    .B_N(net822),
    .Y(_0219_));
 sg13g2_nor3_1 _2744_ (.A(_0871_),
    .B(_0218_),
    .C(_0219_),
    .Y(_0220_));
 sg13g2_nor3_1 _2745_ (.A(net603),
    .B(_0210_),
    .C(_0219_),
    .Y(_0221_));
 sg13g2_nand2_1 _2746_ (.Y(_0222_),
    .A(net839),
    .B(\a[1] ));
 sg13g2_nand2_1 _2747_ (.Y(_0223_),
    .A(net837),
    .B(_0222_));
 sg13g2_o21ai_1 _2748_ (.B1(_0223_),
    .Y(_0224_),
    .A1(_1407_),
    .A2(_0222_));
 sg13g2_o21ai_1 _2749_ (.B1(net822),
    .Y(_0225_),
    .A1(net616),
    .A2(net611));
 sg13g2_nand2b_1 _2750_ (.Y(_0226_),
    .B(net827),
    .A_N(net604));
 sg13g2_nand2_1 _2751_ (.Y(_0227_),
    .A(net606),
    .B(_0223_));
 sg13g2_a22oi_1 _2752_ (.Y(_0228_),
    .B1(_0227_),
    .B2(net827),
    .A2(net622),
    .A1(net737));
 sg13g2_nand2_1 _2753_ (.Y(_0229_),
    .A(_0611_),
    .B(_0228_));
 sg13g2_o21ai_1 _2754_ (.B1(_0226_),
    .Y(_0230_),
    .A1(net827),
    .A2(net837));
 sg13g2_o21ai_1 _2755_ (.B1(_0225_),
    .Y(_0231_),
    .A1(_0621_),
    .A2(_0230_));
 sg13g2_nor4_1 _2756_ (.A(_0220_),
    .B(_0221_),
    .C(_0229_),
    .D(_0231_),
    .Y(_0232_));
 sg13g2_nand2_1 _2757_ (.Y(_0233_),
    .A(_0600_),
    .B(_0198_));
 sg13g2_o21ai_1 _2758_ (.B1(_1568_),
    .Y(uio_out[0]),
    .A1(_0232_),
    .A2(_0233_));
 sg13g2_nand3_1 _2759_ (.B(_1398_),
    .C(_1399_),
    .A(net600),
    .Y(_0234_));
 sg13g2_nand3_1 _2760_ (.B(_1504_),
    .C(_1505_),
    .A(net661),
    .Y(_0235_));
 sg13g2_nand3_1 _2761_ (.B(_1386_),
    .C(_1387_),
    .A(net782),
    .Y(_0236_));
 sg13g2_nand3_1 _2762_ (.B(_1388_),
    .C(_1389_),
    .A(net790),
    .Y(_0237_));
 sg13g2_nand3_1 _2763_ (.B(_0235_),
    .C(_0236_),
    .A(net656),
    .Y(_0238_));
 sg13g2_nand3_1 _2764_ (.B(_0237_),
    .C(_0238_),
    .A(net652),
    .Y(_0239_));
 sg13g2_nand3_1 _2765_ (.B(_1390_),
    .C(_1391_),
    .A(net797),
    .Y(_0240_));
 sg13g2_nand3_1 _2766_ (.B(_1392_),
    .C(_1393_),
    .A(net805),
    .Y(_0241_));
 sg13g2_nand3_1 _2767_ (.B(_0239_),
    .C(_0240_),
    .A(net644),
    .Y(_0242_));
 sg13g2_nand3_1 _2768_ (.B(_0241_),
    .C(_0242_),
    .A(net638),
    .Y(_0243_));
 sg13g2_nand3_1 _2769_ (.B(_1394_),
    .C(_1395_),
    .A(net811),
    .Y(_0244_));
 sg13g2_nand3_1 _2770_ (.B(_1396_),
    .C(_1397_),
    .A(net818),
    .Y(_0245_));
 sg13g2_nand3_1 _2771_ (.B(_0243_),
    .C(_0244_),
    .A(net631),
    .Y(_0246_));
 sg13g2_nand3_1 _2772_ (.B(_0245_),
    .C(_0246_),
    .A(net597),
    .Y(_0247_));
 sg13g2_a21oi_1 _2773_ (.A1(_1280_),
    .A2(_1281_),
    .Y(_0248_),
    .B1(net602));
 sg13g2_a21oi_1 _2774_ (.A1(net734),
    .A2(net615),
    .Y(_0249_),
    .B1(net848));
 sg13g2_a22oi_1 _2775_ (.Y(_0250_),
    .B1(net619),
    .B2(net825),
    .A2(net625),
    .A1(\a[24] ));
 sg13g2_nor2_1 _2776_ (.A(\a[18] ),
    .B(net835),
    .Y(_0251_));
 sg13g2_o21ai_1 _2777_ (.B1(\a[17] ),
    .Y(_0252_),
    .A1(net610),
    .A2(_0251_));
 sg13g2_a21oi_1 _2778_ (.A1(net841),
    .A2(\a[17] ),
    .Y(_0253_),
    .B1(net835));
 sg13g2_o21ai_1 _2779_ (.B1(\a[18] ),
    .Y(_0254_),
    .A1(_1413_),
    .A2(_0253_));
 sg13g2_nand4_1 _2780_ (.B(_0250_),
    .C(_0252_),
    .A(_0249_),
    .Y(_0255_),
    .D(_0254_));
 sg13g2_nor2_1 _2781_ (.A(_0248_),
    .B(_0255_),
    .Y(_0256_));
 sg13g2_nand3_1 _2782_ (.B(_0247_),
    .C(_0256_),
    .A(_0234_),
    .Y(_0257_));
 sg13g2_nor3_1 _2783_ (.A(net639),
    .B(_1545_),
    .C(_1546_),
    .Y(_0258_));
 sg13g2_nand3_1 _2784_ (.B(_1543_),
    .C(_1544_),
    .A(net803),
    .Y(_0259_));
 sg13g2_a21o_1 _2785_ (.A2(_1539_),
    .A1(net784),
    .B1(net789),
    .X(_0260_));
 sg13g2_o21ai_1 _2786_ (.B1(net789),
    .Y(_0261_),
    .A1(_1540_),
    .A2(_1541_));
 sg13g2_nand3_1 _2787_ (.B(_0260_),
    .C(_0261_),
    .A(net649),
    .Y(_0262_));
 sg13g2_nand3_1 _2788_ (.B(_1538_),
    .C(_1542_),
    .A(net798),
    .Y(_0263_));
 sg13g2_nand3_1 _2789_ (.B(_0262_),
    .C(_0263_),
    .A(net645),
    .Y(_0264_));
 sg13g2_a21oi_1 _2790_ (.A1(_0259_),
    .A2(_0264_),
    .Y(_0265_),
    .B1(net812));
 sg13g2_a21oi_1 _2791_ (.A1(_1034_),
    .A2(_1035_),
    .Y(_0266_),
    .B1(net602));
 sg13g2_a21oi_1 _2792_ (.A1(\a[28] ),
    .A2(net624),
    .Y(_0267_),
    .B1(_0611_));
 sg13g2_a22oi_1 _2793_ (.Y(_0268_),
    .B1(net614),
    .B2(net717),
    .A2(net619),
    .A1(\a[12] ));
 sg13g2_and2_1 _2794_ (.A(net842),
    .B(\a[26] ),
    .X(_0269_));
 sg13g2_nor2_1 _2795_ (.A(net834),
    .B(_0269_),
    .Y(_0270_));
 sg13g2_a21oi_1 _2796_ (.A1(\a[25] ),
    .A2(_0269_),
    .Y(_0271_),
    .B1(net834));
 sg13g2_o21ai_1 _2797_ (.B1(_0271_),
    .Y(_0272_),
    .A1(\a[25] ),
    .A2(\a[26] ));
 sg13g2_and2_1 _2798_ (.A(_1406_),
    .B(_0269_),
    .X(_0273_));
 sg13g2_o21ai_1 _2799_ (.B1(\a[25] ),
    .Y(_0274_),
    .A1(net610),
    .A2(_0273_));
 sg13g2_nand4_1 _2800_ (.B(_0268_),
    .C(_0272_),
    .A(_0267_),
    .Y(_0275_),
    .D(_0274_));
 sg13g2_nor2_1 _2801_ (.A(_0266_),
    .B(_0275_),
    .Y(_0276_));
 sg13g2_nor3_1 _2802_ (.A(net649),
    .B(_1550_),
    .C(_1551_),
    .Y(_0277_));
 sg13g2_a21oi_1 _2803_ (.A1(_0260_),
    .A2(_0261_),
    .Y(_0278_),
    .B1(net798));
 sg13g2_nor3_1 _2804_ (.A(net803),
    .B(_0277_),
    .C(_0278_),
    .Y(_0279_));
 sg13g2_a21oi_1 _2805_ (.A1(net806),
    .A2(_1553_),
    .Y(_0280_),
    .B1(_0279_));
 sg13g2_mux2_1 _2806_ (.A0(_1554_),
    .A1(_0280_),
    .S(net636),
    .X(_0281_));
 sg13g2_mux2_1 _2807_ (.A0(_1555_),
    .A1(_0281_),
    .S(net632),
    .X(_0282_));
 sg13g2_o21ai_1 _2808_ (.B1(_0276_),
    .Y(_0283_),
    .A1(_1371_),
    .A2(_0282_));
 sg13g2_a21oi_1 _2809_ (.A1(net601),
    .A2(_1556_),
    .Y(_0284_),
    .B1(_0283_));
 sg13g2_nand2_1 _2810_ (.Y(_0285_),
    .A(net843),
    .B(_0257_));
 sg13g2_nand3_1 _2811_ (.B(_0090_),
    .C(_0091_),
    .A(net599),
    .Y(_0286_));
 sg13g2_nand3_1 _2812_ (.B(_1355_),
    .C(_1356_),
    .A(net661),
    .Y(_0287_));
 sg13g2_nand3_1 _2813_ (.B(_1675_),
    .C(_1676_),
    .A(net782),
    .Y(_0288_));
 sg13g2_nand3_1 _2814_ (.B(_1677_),
    .C(_0064_),
    .A(net789),
    .Y(_0289_));
 sg13g2_nand3_1 _2815_ (.B(_0287_),
    .C(_0288_),
    .A(net656),
    .Y(_0290_));
 sg13g2_nand3_1 _2816_ (.B(_0289_),
    .C(_0290_),
    .A(net652),
    .Y(_0291_));
 sg13g2_nand3_1 _2817_ (.B(_0065_),
    .C(_0066_),
    .A(net798),
    .Y(_0292_));
 sg13g2_nand3_1 _2818_ (.B(_0067_),
    .C(_0068_),
    .A(net803),
    .Y(_0293_));
 sg13g2_nand3_1 _2819_ (.B(_0291_),
    .C(_0292_),
    .A(net645),
    .Y(_0294_));
 sg13g2_nand3_1 _2820_ (.B(_0293_),
    .C(_0294_),
    .A(net636),
    .Y(_0295_));
 sg13g2_nand3_1 _2821_ (.B(_0069_),
    .C(_0070_),
    .A(net809),
    .Y(_0296_));
 sg13g2_nand3_1 _2822_ (.B(_0071_),
    .C(_0072_),
    .A(net815),
    .Y(_0297_));
 sg13g2_nand3_1 _2823_ (.B(_0295_),
    .C(_0296_),
    .A(net632),
    .Y(_0298_));
 sg13g2_nand3_1 _2824_ (.B(_0297_),
    .C(_0298_),
    .A(net594),
    .Y(_0299_));
 sg13g2_a21oi_1 _2825_ (.A1(\a[4] ),
    .A2(net617),
    .Y(_0300_),
    .B1(_0611_));
 sg13g2_a22oi_1 _2826_ (.Y(_0301_),
    .B1(net613),
    .B2(net767),
    .A2(net622),
    .A1(\a[20] ));
 sg13g2_and2_1 _2827_ (.A(\a[10] ),
    .B(net604),
    .X(_0302_));
 sg13g2_o21ai_1 _2828_ (.B1(\a[9] ),
    .Y(_0303_),
    .A1(net609),
    .A2(_0302_));
 sg13g2_a21oi_1 _2829_ (.A1(net839),
    .A2(\a[10] ),
    .Y(_0304_),
    .B1(net832));
 sg13g2_or2_1 _2830_ (.X(_0305_),
    .B(\a[10] ),
    .A(\a[9] ));
 sg13g2_o21ai_1 _2831_ (.B1(_0305_),
    .Y(_0306_),
    .A1(_0185_),
    .A2(_0304_));
 sg13g2_nand4_1 _2832_ (.B(_0301_),
    .C(_0303_),
    .A(_0300_),
    .Y(_0307_),
    .D(_0306_));
 sg13g2_nor3_1 _2833_ (.A(net659),
    .B(net786),
    .C(_0189_),
    .Y(_0308_));
 sg13g2_a21oi_1 _2834_ (.A1(net786),
    .A2(_0191_),
    .Y(_0309_),
    .B1(_0308_));
 sg13g2_nand2_1 _2835_ (.Y(_0310_),
    .A(net793),
    .B(_0192_));
 sg13g2_o21ai_1 _2836_ (.B1(_0310_),
    .Y(_0311_),
    .A1(net793),
    .A2(_0309_));
 sg13g2_mux2_1 _2837_ (.A0(_0193_),
    .A1(_0311_),
    .S(net640),
    .X(_0312_));
 sg13g2_mux2_1 _2838_ (.A0(_0194_),
    .A1(_0312_),
    .S(net633),
    .X(_0313_));
 sg13g2_mux2_1 _2839_ (.A0(_0195_),
    .A1(_0313_),
    .S(net628),
    .X(_0314_));
 sg13g2_a221oi_1 _2840_ (.B2(net589),
    .C1(_0307_),
    .B1(_0314_),
    .A1(net591),
    .Y(_0315_),
    .A2(_0196_));
 sg13g2_nand3_1 _2841_ (.B(_0299_),
    .C(_0315_),
    .A(_0286_),
    .Y(_0316_));
 sg13g2_nand3b_1 _2842_ (.B(_0216_),
    .C(net816),
    .Y(_0317_),
    .A_N(_0207_));
 sg13g2_nor2_1 _2843_ (.A(net640),
    .B(_0204_),
    .Y(_0318_));
 sg13g2_nand2_1 _2844_ (.Y(_0319_),
    .A(_0214_),
    .B(_0318_));
 sg13g2_nor2_1 _2845_ (.A(net654),
    .B(_0201_),
    .Y(_0320_));
 sg13g2_nand2_1 _2846_ (.Y(_0321_),
    .A(_0212_),
    .B(_0320_));
 sg13g2_a21oi_1 _2847_ (.A1(_0097_),
    .A2(_0098_),
    .Y(_0322_),
    .B1(net781));
 sg13g2_nor3_1 _2848_ (.A(net659),
    .B(_0200_),
    .C(_0211_),
    .Y(_0323_));
 sg13g2_o21ai_1 _2849_ (.B1(net655),
    .Y(_0324_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_a21oi_1 _2850_ (.A1(_0321_),
    .A2(_0324_),
    .Y(_0325_),
    .B1(net795));
 sg13g2_nor3_1 _2851_ (.A(net646),
    .B(_0203_),
    .C(_0213_),
    .Y(_0326_));
 sg13g2_o21ai_1 _2852_ (.B1(net640),
    .Y(_0327_),
    .A1(_0325_),
    .A2(_0326_));
 sg13g2_a21oi_1 _2853_ (.A1(_0319_),
    .A2(_0327_),
    .Y(_0328_),
    .B1(net808));
 sg13g2_nand2b_1 _2854_ (.Y(_0329_),
    .B(net808),
    .A_N(_0206_));
 sg13g2_nor2_1 _2855_ (.A(_0215_),
    .B(_0329_),
    .Y(_0330_));
 sg13g2_o21ai_1 _2856_ (.B1(net626),
    .Y(_0331_),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_a21oi_1 _2857_ (.A1(_0317_),
    .A2(_0331_),
    .Y(_0332_),
    .B1(net822));
 sg13g2_nand2b_1 _2858_ (.Y(_0333_),
    .B(net822),
    .A_N(_0209_));
 sg13g2_o21ai_1 _2859_ (.B1(_0870_),
    .Y(_0334_),
    .A1(_0217_),
    .A2(_0333_));
 sg13g2_mux2_1 _2860_ (.A0(_0166_),
    .A1(_0200_),
    .S(net780),
    .X(_0335_));
 sg13g2_nor2_1 _2861_ (.A(net786),
    .B(_0335_),
    .Y(_0336_));
 sg13g2_nor2_1 _2862_ (.A(_0320_),
    .B(_0336_),
    .Y(_0337_));
 sg13g2_mux2_1 _2863_ (.A0(_0203_),
    .A1(_0337_),
    .S(net647),
    .X(_0338_));
 sg13g2_nor2_1 _2864_ (.A(net802),
    .B(_0338_),
    .Y(_0339_));
 sg13g2_nor2_1 _2865_ (.A(_0318_),
    .B(_0339_),
    .Y(_0340_));
 sg13g2_o21ai_1 _2866_ (.B1(_0329_),
    .Y(_0341_),
    .A1(net808),
    .A2(_0340_));
 sg13g2_nand2_1 _2867_ (.Y(_0342_),
    .A(net626),
    .B(_0341_));
 sg13g2_o21ai_1 _2868_ (.B1(_0342_),
    .Y(_0343_),
    .A1(net627),
    .A2(_0207_));
 sg13g2_inv_1 _2869_ (.Y(_0344_),
    .A(_0343_));
 sg13g2_nor2_1 _2870_ (.A(\a[2] ),
    .B(net832),
    .Y(_0345_));
 sg13g2_o21ai_1 _2871_ (.B1(\a[1] ),
    .Y(_0346_),
    .A1(net608),
    .A2(_0345_));
 sg13g2_a221oi_1 _2872_ (.B2(net816),
    .C1(net845),
    .B1(net611),
    .A1(net830),
    .Y(_0347_),
    .A2(net621));
 sg13g2_a22oi_1 _2873_ (.Y(_0348_),
    .B1(_0224_),
    .B2(\a[2] ),
    .A2(net616),
    .A1(net828));
 sg13g2_nand3_1 _2874_ (.B(_0347_),
    .C(_0348_),
    .A(_0346_),
    .Y(_0349_));
 sg13g2_a221oi_1 _2875_ (.B2(net589),
    .C1(_0349_),
    .B1(_0344_),
    .A1(net591),
    .Y(_0350_),
    .A2(_0209_));
 sg13g2_o21ai_1 _2876_ (.B1(_0350_),
    .Y(_0351_),
    .A1(_0332_),
    .A2(_0334_));
 sg13g2_nand3_1 _2877_ (.B(_0316_),
    .C(_0351_),
    .A(_0600_),
    .Y(_0352_));
 sg13g2_o21ai_1 _2878_ (.B1(_0352_),
    .Y(uio_out[1]),
    .A1(_0284_),
    .A2(_0285_));
 sg13g2_nand3_1 _2879_ (.B(_0235_),
    .C(_0236_),
    .A(net790),
    .Y(_0353_));
 sg13g2_nand3_1 _2880_ (.B(_1506_),
    .C(_1507_),
    .A(net656),
    .Y(_0354_));
 sg13g2_nand3_1 _2881_ (.B(_0353_),
    .C(_0354_),
    .A(net651),
    .Y(_0355_));
 sg13g2_nand3_1 _2882_ (.B(_0237_),
    .C(_0238_),
    .A(net796),
    .Y(_0356_));
 sg13g2_nand3_1 _2883_ (.B(_0239_),
    .C(_0240_),
    .A(net805),
    .Y(_0357_));
 sg13g2_nand3_1 _2884_ (.B(_0355_),
    .C(_0356_),
    .A(net643),
    .Y(_0358_));
 sg13g2_nand3_1 _2885_ (.B(_0357_),
    .C(_0358_),
    .A(net637),
    .Y(_0359_));
 sg13g2_nand3_1 _2886_ (.B(_0241_),
    .C(_0242_),
    .A(net811),
    .Y(_0360_));
 sg13g2_nand3_1 _2887_ (.B(_0243_),
    .C(_0244_),
    .A(net819),
    .Y(_0361_));
 sg13g2_nand3_1 _2888_ (.B(_0359_),
    .C(_0360_),
    .A(net631),
    .Y(_0362_));
 sg13g2_nand3_1 _2889_ (.B(_0361_),
    .C(_0362_),
    .A(net596),
    .Y(_0363_));
 sg13g2_nand3_1 _2890_ (.B(_0245_),
    .C(_0246_),
    .A(net600),
    .Y(_0364_));
 sg13g2_a21oi_1 _2891_ (.A1(_1226_),
    .A2(_1227_),
    .Y(_0365_),
    .B1(net602));
 sg13g2_a22oi_1 _2892_ (.Y(_0366_),
    .B1(net620),
    .B2(net767),
    .A2(net623),
    .A1(net717));
 sg13g2_a21oi_1 _2893_ (.A1(net730),
    .A2(net614),
    .Y(_0367_),
    .B1(net849));
 sg13g2_and2_1 _2894_ (.A(net841),
    .B(\a[19] ),
    .X(_0368_));
 sg13g2_nor2_1 _2895_ (.A(net834),
    .B(_0368_),
    .Y(_0369_));
 sg13g2_a21oi_1 _2896_ (.A1(\a[18] ),
    .A2(_0368_),
    .Y(_0370_),
    .B1(net834));
 sg13g2_o21ai_1 _2897_ (.B1(_0370_),
    .Y(_0371_),
    .A1(\a[18] ),
    .A2(\a[19] ));
 sg13g2_and2_1 _2898_ (.A(_1406_),
    .B(_0368_),
    .X(_0372_));
 sg13g2_o21ai_1 _2899_ (.B1(\a[18] ),
    .Y(_0373_),
    .A1(net610),
    .A2(_0372_));
 sg13g2_nand4_1 _2900_ (.B(_0367_),
    .C(_0371_),
    .A(_0366_),
    .Y(_0374_),
    .D(_0373_));
 sg13g2_nor2_1 _2901_ (.A(_0365_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_nand3_1 _2902_ (.B(_0364_),
    .C(_0375_),
    .A(_0363_),
    .Y(_0376_));
 sg13g2_nand3_1 _2903_ (.B(_0262_),
    .C(_0263_),
    .A(net803),
    .Y(_0377_));
 sg13g2_nand3_1 _2904_ (.B(net789),
    .C(_1539_),
    .A(net784),
    .Y(_0378_));
 sg13g2_and2_1 _2905_ (.A(net649),
    .B(_0378_),
    .X(_0379_));
 sg13g2_a21oi_1 _2906_ (.A1(_0260_),
    .A2(_0261_),
    .Y(_0380_),
    .B1(net649));
 sg13g2_o21ai_1 _2907_ (.B1(net645),
    .Y(_0381_),
    .A1(_0379_),
    .A2(_0380_));
 sg13g2_nand3_1 _2908_ (.B(_0377_),
    .C(_0381_),
    .A(net636),
    .Y(_0382_));
 sg13g2_nand3_1 _2909_ (.B(_0259_),
    .C(_0264_),
    .A(net812),
    .Y(_0383_));
 sg13g2_nand2_1 _2910_ (.Y(_0384_),
    .A(_0382_),
    .B(_0383_));
 sg13g2_nor3_1 _2911_ (.A(net632),
    .B(_0258_),
    .C(_0265_),
    .Y(_0385_));
 sg13g2_a21oi_1 _2912_ (.A1(net632),
    .A2(_0384_),
    .Y(_0386_),
    .B1(_0385_));
 sg13g2_nor2_1 _2913_ (.A(_1371_),
    .B(_0386_),
    .Y(_0387_));
 sg13g2_nor2_1 _2914_ (.A(_0873_),
    .B(_0282_),
    .Y(_0388_));
 sg13g2_a22oi_1 _2915_ (.Y(_0389_),
    .B1(net620),
    .B2(net748),
    .A2(net623),
    .A1(\ayayayayayaya.b[29] ));
 sg13g2_inv_1 _2916_ (.Y(_0390_),
    .A(_0389_));
 sg13g2_nor2_1 _2917_ (.A(\a[27] ),
    .B(net834),
    .Y(_0391_));
 sg13g2_o21ai_1 _2918_ (.B1(\a[26] ),
    .Y(_0392_),
    .A1(net610),
    .A2(_0391_));
 sg13g2_o21ai_1 _2919_ (.B1(\a[27] ),
    .Y(_0393_),
    .A1(_0270_),
    .A2(_0273_));
 sg13g2_a221oi_1 _2920_ (.B2(_1071_),
    .C1(_0390_),
    .B1(_1423_),
    .A1(net716),
    .Y(_0394_),
    .A2(net615));
 sg13g2_nand4_1 _2921_ (.B(_0392_),
    .C(_0393_),
    .A(net848),
    .Y(_0395_),
    .D(_0394_));
 sg13g2_nor3_1 _2922_ (.A(_0387_),
    .B(_0388_),
    .C(_0395_),
    .Y(_0396_));
 sg13g2_nand2_1 _2923_ (.Y(_0397_),
    .A(net843),
    .B(_0376_));
 sg13g2_nand3_1 _2924_ (.B(_0297_),
    .C(_0298_),
    .A(net599),
    .Y(_0398_));
 sg13g2_nand3_1 _2925_ (.B(_0287_),
    .C(_0288_),
    .A(net790),
    .Y(_0399_));
 sg13g2_nand3_1 _2926_ (.B(_1357_),
    .C(_1358_),
    .A(net656),
    .Y(_0400_));
 sg13g2_nand3_1 _2927_ (.B(_0399_),
    .C(_0400_),
    .A(net652),
    .Y(_0401_));
 sg13g2_nand3_1 _2928_ (.B(_0289_),
    .C(_0290_),
    .A(net796),
    .Y(_0402_));
 sg13g2_nand3_1 _2929_ (.B(_0291_),
    .C(_0292_),
    .A(net803),
    .Y(_0403_));
 sg13g2_nand3_1 _2930_ (.B(_0401_),
    .C(_0402_),
    .A(net643),
    .Y(_0404_));
 sg13g2_nand3_1 _2931_ (.B(_0403_),
    .C(_0404_),
    .A(net636),
    .Y(_0405_));
 sg13g2_nand3_1 _2932_ (.B(_0293_),
    .C(_0294_),
    .A(net812),
    .Y(_0406_));
 sg13g2_nand3_1 _2933_ (.B(_0295_),
    .C(_0296_),
    .A(net815),
    .Y(_0407_));
 sg13g2_nand3_1 _2934_ (.B(_0405_),
    .C(_0406_),
    .A(net632),
    .Y(_0408_));
 sg13g2_and2_1 _2935_ (.A(_0407_),
    .B(_0408_),
    .X(_0409_));
 sg13g2_nand3_1 _2936_ (.B(_0407_),
    .C(_0408_),
    .A(net593),
    .Y(_0410_));
 sg13g2_nand2_1 _2937_ (.Y(_0411_),
    .A(net762),
    .B(net611));
 sg13g2_o21ai_1 _2938_ (.B1(\a[11] ),
    .Y(_0412_),
    .A1(_0302_),
    .A2(_0304_));
 sg13g2_nor2_1 _2939_ (.A(\a[11] ),
    .B(net833),
    .Y(_0413_));
 sg13g2_o21ai_1 _2940_ (.B1(\a[10] ),
    .Y(_0414_),
    .A1(net608),
    .A2(_0413_));
 sg13g2_nand4_1 _2941_ (.B(_0411_),
    .C(_0412_),
    .A(net845),
    .Y(_0415_),
    .D(_0414_));
 sg13g2_a221oi_1 _2942_ (.B2(net788),
    .C1(_0415_),
    .B1(net618),
    .A1(net724),
    .Y(_0416_),
    .A2(net622));
 sg13g2_nor2_1 _2943_ (.A(net640),
    .B(_0311_),
    .Y(_0417_));
 sg13g2_nor3_1 _2944_ (.A(net659),
    .B(net654),
    .C(_0189_),
    .Y(_0418_));
 sg13g2_nor2_1 _2945_ (.A(net646),
    .B(_0309_),
    .Y(_0419_));
 sg13g2_a21oi_1 _2946_ (.A1(net648),
    .A2(_0418_),
    .Y(_0420_),
    .B1(_0419_));
 sg13g2_a21oi_1 _2947_ (.A1(net642),
    .A2(_0420_),
    .Y(_0421_),
    .B1(_0417_));
 sg13g2_mux2_1 _2948_ (.A0(_0312_),
    .A1(_0421_),
    .S(net633),
    .X(_0422_));
 sg13g2_mux2_1 _2949_ (.A0(_0313_),
    .A1(_0422_),
    .S(net627),
    .X(_0423_));
 sg13g2_a22oi_1 _2950_ (.Y(_0424_),
    .B1(_0423_),
    .B2(net590),
    .A2(_0314_),
    .A1(net592));
 sg13g2_nand4_1 _2951_ (.B(_0410_),
    .C(_0416_),
    .A(_0398_),
    .Y(_0425_),
    .D(_0424_));
 sg13g2_o21ai_1 _2952_ (.B1(net786),
    .Y(_0426_),
    .A1(_0322_),
    .A2(_0323_));
 sg13g2_nand3_1 _2953_ (.B(_0099_),
    .C(_0100_),
    .A(net654),
    .Y(_0427_));
 sg13g2_nand3_1 _2954_ (.B(_0426_),
    .C(_0427_),
    .A(net646),
    .Y(_0428_));
 sg13g2_nand3_1 _2955_ (.B(_0321_),
    .C(_0324_),
    .A(net793),
    .Y(_0429_));
 sg13g2_o21ai_1 _2956_ (.B1(net802),
    .Y(_0430_),
    .A1(_0325_),
    .A2(_0326_));
 sg13g2_nand3_1 _2957_ (.B(_0428_),
    .C(_0429_),
    .A(net641),
    .Y(_0431_));
 sg13g2_nand3_1 _2958_ (.B(_0430_),
    .C(_0431_),
    .A(net634),
    .Y(_0432_));
 sg13g2_nand3_1 _2959_ (.B(_0319_),
    .C(_0327_),
    .A(net808),
    .Y(_0433_));
 sg13g2_o21ai_1 _2960_ (.B1(net816),
    .Y(_0434_),
    .A1(_0328_),
    .A2(_0330_));
 sg13g2_nand3_1 _2961_ (.B(_0432_),
    .C(_0433_),
    .A(net627),
    .Y(_0435_));
 sg13g2_and2_1 _2962_ (.A(_0434_),
    .B(_0435_),
    .X(_0436_));
 sg13g2_nand3_1 _2963_ (.B(_0434_),
    .C(_0435_),
    .A(net593),
    .Y(_0437_));
 sg13g2_nand3_1 _2964_ (.B(_0317_),
    .C(_0331_),
    .A(net598),
    .Y(_0438_));
 sg13g2_mux2_1 _2965_ (.A0(_0167_),
    .A1(_0335_),
    .S(net787),
    .X(_0439_));
 sg13g2_mux2_1 _2966_ (.A0(_0337_),
    .A1(_0439_),
    .S(net647),
    .X(_0440_));
 sg13g2_mux2_1 _2967_ (.A0(_0338_),
    .A1(_0440_),
    .S(net641),
    .X(_0441_));
 sg13g2_mux2_1 _2968_ (.A0(_0340_),
    .A1(_0441_),
    .S(net634),
    .X(_0442_));
 sg13g2_nor2_1 _2969_ (.A(net816),
    .B(_0442_),
    .Y(_0443_));
 sg13g2_a21oi_1 _2970_ (.A1(net816),
    .A2(_0341_),
    .Y(_0444_),
    .B1(_0443_));
 sg13g2_a21o_1 _2971_ (.A2(net617),
    .A1(net817),
    .B1(net845),
    .X(_0445_));
 sg13g2_a221oi_1 _2972_ (.B2(net808),
    .C1(_0445_),
    .B1(net611),
    .A1(net734),
    .Y(_0446_),
    .A2(net621));
 sg13g2_and2_1 _2973_ (.A(\a[3] ),
    .B(net604),
    .X(_0447_));
 sg13g2_o21ai_1 _2974_ (.B1(\a[2] ),
    .Y(_0448_),
    .A1(net608),
    .A2(_0447_));
 sg13g2_a21oi_1 _2975_ (.A1(net839),
    .A2(\a[3] ),
    .Y(_0449_),
    .B1(net832));
 sg13g2_or2_1 _2976_ (.X(_0450_),
    .B(\a[3] ),
    .A(\a[2] ));
 sg13g2_o21ai_1 _2977_ (.B1(_0450_),
    .Y(_0451_),
    .A1(_0345_),
    .A2(_0449_));
 sg13g2_nand3_1 _2978_ (.B(_0448_),
    .C(_0451_),
    .A(_0446_),
    .Y(_0452_));
 sg13g2_a221oi_1 _2979_ (.B2(net589),
    .C1(_0452_),
    .B1(_0444_),
    .A1(net591),
    .Y(_0453_),
    .A2(_0344_));
 sg13g2_nand3_1 _2980_ (.B(_0438_),
    .C(_0453_),
    .A(_0437_),
    .Y(_0454_));
 sg13g2_nand3_1 _2981_ (.B(_0425_),
    .C(_0454_),
    .A(_0600_),
    .Y(_0455_));
 sg13g2_o21ai_1 _2982_ (.B1(_0455_),
    .Y(uio_out[2]),
    .A1(_0396_),
    .A2(_0397_));
 sg13g2_nand3_1 _2983_ (.B(_1508_),
    .C(_1509_),
    .A(net651),
    .Y(_0456_));
 sg13g2_nand3_1 _2984_ (.B(_0353_),
    .C(_0354_),
    .A(net796),
    .Y(_0457_));
 sg13g2_nand3_1 _2985_ (.B(_0355_),
    .C(_0356_),
    .A(net805),
    .Y(_0458_));
 sg13g2_nand3_1 _2986_ (.B(_0456_),
    .C(_0457_),
    .A(net643),
    .Y(_0459_));
 sg13g2_nand3_1 _2987_ (.B(_0458_),
    .C(_0459_),
    .A(net637),
    .Y(_0460_));
 sg13g2_nand3_1 _2988_ (.B(_0357_),
    .C(_0358_),
    .A(net811),
    .Y(_0461_));
 sg13g2_nand3_1 _2989_ (.B(_0359_),
    .C(_0360_),
    .A(net819),
    .Y(_0462_));
 sg13g2_nand3_1 _2990_ (.B(_0460_),
    .C(_0461_),
    .A(net631),
    .Y(_0463_));
 sg13g2_nand3_1 _2991_ (.B(_0462_),
    .C(_0463_),
    .A(net595),
    .Y(_0464_));
 sg13g2_a21oi_1 _2992_ (.A1(_1177_),
    .A2(_1178_),
    .Y(_0465_),
    .B1(net602));
 sg13g2_o21ai_1 _2993_ (.B1(\a[20] ),
    .Y(_0466_),
    .A1(_0369_),
    .A2(_0372_));
 sg13g2_o21ai_1 _2994_ (.B1(net606),
    .Y(_0467_),
    .A1(\a[20] ),
    .A2(net832));
 sg13g2_a22oi_1 _2995_ (.Y(_0468_),
    .B1(net614),
    .B2(net728),
    .A2(net624),
    .A1(\a[25] ));
 sg13g2_a22oi_1 _2996_ (.Y(_0469_),
    .B1(_0467_),
    .B2(\a[19] ),
    .A2(net617),
    .A1(\a[9] ));
 sg13g2_nand4_1 _2997_ (.B(_0466_),
    .C(_0468_),
    .A(_0611_),
    .Y(_0470_),
    .D(_0469_));
 sg13g2_nor2_1 _2998_ (.A(_0465_),
    .B(_0470_),
    .Y(_0471_));
 sg13g2_nand3_1 _2999_ (.B(_0361_),
    .C(_0362_),
    .A(net600),
    .Y(_0472_));
 sg13g2_nand3_1 _3000_ (.B(_0471_),
    .C(_0472_),
    .A(_0464_),
    .Y(_0473_));
 sg13g2_o21ai_1 _3001_ (.B1(net645),
    .Y(_0474_),
    .A1(net650),
    .A2(_0378_));
 sg13g2_o21ai_1 _3002_ (.B1(net806),
    .Y(_0475_),
    .A1(_0379_),
    .A2(_0380_));
 sg13g2_nand3_1 _3003_ (.B(_0474_),
    .C(_0475_),
    .A(net636),
    .Y(_0476_));
 sg13g2_nand3_1 _3004_ (.B(_0377_),
    .C(_0381_),
    .A(net812),
    .Y(_0477_));
 sg13g2_nand2_1 _3005_ (.Y(_0478_),
    .A(_0476_),
    .B(_0477_));
 sg13g2_mux2_1 _3006_ (.A0(_0384_),
    .A1(_0478_),
    .S(net632),
    .X(_0479_));
 sg13g2_nand2_1 _3007_ (.Y(_0480_),
    .A(\ayayayayayaya.b[27] ),
    .B(net614));
 sg13g2_a22oi_1 _3008_ (.Y(_0481_),
    .B1(net619),
    .B2(\a[13] ),
    .A2(net625),
    .A1(\a[29] ));
 sg13g2_nand2_1 _3009_ (.Y(_0482_),
    .A(net841),
    .B(\a[28] ));
 sg13g2_a21o_1 _3010_ (.A2(_0482_),
    .A1(net837),
    .B1(_0391_),
    .X(_0483_));
 sg13g2_o21ai_1 _3011_ (.B1(_0483_),
    .Y(_0484_),
    .A1(\a[27] ),
    .A2(\a[28] ));
 sg13g2_o21ai_1 _3012_ (.B1(net607),
    .Y(_0485_),
    .A1(_1407_),
    .A2(_0482_));
 sg13g2_nand4_1 _3013_ (.B(_0480_),
    .C(_0481_),
    .A(net848),
    .Y(_0486_),
    .D(_0484_));
 sg13g2_a221oi_1 _3014_ (.B2(\a[27] ),
    .C1(_0486_),
    .B1(_0485_),
    .A1(_1111_),
    .Y(_0487_),
    .A2(_1423_));
 sg13g2_o21ai_1 _3015_ (.B1(_0487_),
    .Y(_0488_),
    .A1(_0873_),
    .A2(_0386_));
 sg13g2_a21oi_1 _3016_ (.A1(net596),
    .A2(_0479_),
    .Y(_0489_),
    .B1(_0488_));
 sg13g2_nand2_1 _3017_ (.Y(_0490_),
    .A(net844),
    .B(_0473_));
 sg13g2_nand3_1 _3018_ (.B(_1359_),
    .C(_1360_),
    .A(net651),
    .Y(_0491_));
 sg13g2_nand3_1 _3019_ (.B(_0399_),
    .C(_0400_),
    .A(net796),
    .Y(_0492_));
 sg13g2_nand3_1 _3020_ (.B(_0401_),
    .C(_0402_),
    .A(net804),
    .Y(_0493_));
 sg13g2_nand3_1 _3021_ (.B(_0491_),
    .C(_0492_),
    .A(net644),
    .Y(_0494_));
 sg13g2_nand3_1 _3022_ (.B(_0493_),
    .C(_0494_),
    .A(net637),
    .Y(_0495_));
 sg13g2_nand3_1 _3023_ (.B(_0403_),
    .C(_0404_),
    .A(net812),
    .Y(_0496_));
 sg13g2_a21oi_1 _3024_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0497_),
    .B1(net820));
 sg13g2_a21oi_1 _3025_ (.A1(_0405_),
    .A2(_0406_),
    .Y(_0498_),
    .B1(net632));
 sg13g2_or2_1 _3026_ (.X(_0499_),
    .B(_0498_),
    .A(_0497_));
 sg13g2_nand2_1 _3027_ (.Y(_0500_),
    .A(\a[5] ),
    .B(net616));
 sg13g2_nand2_1 _3028_ (.Y(_0501_),
    .A(net845),
    .B(_0500_));
 sg13g2_a221oi_1 _3029_ (.B2(net754),
    .C1(_0501_),
    .B1(net611),
    .A1(\a[21] ),
    .Y(_0502_),
    .A2(net621));
 sg13g2_and2_1 _3030_ (.A(\a[12] ),
    .B(net605),
    .X(_0503_));
 sg13g2_o21ai_1 _3031_ (.B1(\a[11] ),
    .Y(_0504_),
    .A1(net609),
    .A2(_0503_));
 sg13g2_a21oi_1 _3032_ (.A1(net839),
    .A2(\a[12] ),
    .Y(_0505_),
    .B1(net833));
 sg13g2_or2_1 _3033_ (.X(_0506_),
    .B(\a[12] ),
    .A(\a[11] ));
 sg13g2_o21ai_1 _3034_ (.B1(_0506_),
    .Y(_0507_),
    .A1(_0413_),
    .A2(_0505_));
 sg13g2_a21oi_1 _3035_ (.A1(net794),
    .A2(_0418_),
    .Y(_0508_),
    .B1(net800));
 sg13g2_a21oi_1 _3036_ (.A1(net800),
    .A2(_0420_),
    .Y(_0509_),
    .B1(_0508_));
 sg13g2_mux2_1 _3037_ (.A0(_0421_),
    .A1(_0509_),
    .S(net635),
    .X(_0510_));
 sg13g2_mux2_1 _3038_ (.A0(_0422_),
    .A1(_0510_),
    .S(net629),
    .X(_0511_));
 sg13g2_a22oi_1 _3039_ (.Y(_0512_),
    .B1(_0511_),
    .B2(net590),
    .A2(_0423_),
    .A1(net592));
 sg13g2_nand4_1 _3040_ (.B(_0504_),
    .C(_0507_),
    .A(_0502_),
    .Y(_0513_),
    .D(_0512_));
 sg13g2_a221oi_1 _3041_ (.B2(net593),
    .C1(_0513_),
    .B1(_0499_),
    .A1(net599),
    .Y(_0514_),
    .A2(_0409_));
 sg13g2_nand3_1 _3042_ (.B(_0101_),
    .C(_0102_),
    .A(net646),
    .Y(_0515_));
 sg13g2_nand3_1 _3043_ (.B(_0426_),
    .C(_0427_),
    .A(net794),
    .Y(_0516_));
 sg13g2_nand3_1 _3044_ (.B(_0428_),
    .C(_0429_),
    .A(net800),
    .Y(_0517_));
 sg13g2_nand3_1 _3045_ (.B(_0515_),
    .C(_0516_),
    .A(net641),
    .Y(_0518_));
 sg13g2_nand3_1 _3046_ (.B(_0517_),
    .C(_0518_),
    .A(net634),
    .Y(_0519_));
 sg13g2_nand3_1 _3047_ (.B(_0430_),
    .C(_0431_),
    .A(net808),
    .Y(_0520_));
 sg13g2_a21oi_1 _3048_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0521_),
    .B1(net814));
 sg13g2_a21oi_1 _3049_ (.A1(_0432_),
    .A2(_0433_),
    .Y(_0522_),
    .B1(net626));
 sg13g2_or2_1 _3050_ (.X(_0523_),
    .B(_0522_),
    .A(_0521_));
 sg13g2_a21o_1 _3051_ (.A2(net616),
    .A1(\a[1] ),
    .B1(net845),
    .X(_0524_));
 sg13g2_a221oi_1 _3052_ (.B2(net802),
    .C1(_0524_),
    .B1(net611),
    .A1(\a[17] ),
    .Y(_0525_),
    .A2(net621));
 sg13g2_o21ai_1 _3053_ (.B1(\a[4] ),
    .Y(_0526_),
    .A1(_0447_),
    .A2(_0449_));
 sg13g2_nor2_1 _3054_ (.A(\a[4] ),
    .B(net832),
    .Y(_0527_));
 sg13g2_o21ai_1 _3055_ (.B1(\a[3] ),
    .Y(_0528_),
    .A1(net608),
    .A2(_0527_));
 sg13g2_mux2_1 _3056_ (.A0(_0168_),
    .A1(_0439_),
    .S(net793),
    .X(_0529_));
 sg13g2_mux2_1 _3057_ (.A0(_0440_),
    .A1(_0529_),
    .S(net641),
    .X(_0530_));
 sg13g2_mux2_1 _3058_ (.A0(_0441_),
    .A1(_0530_),
    .S(net634),
    .X(_0531_));
 sg13g2_mux2_1 _3059_ (.A0(_0442_),
    .A1(_0531_),
    .S(net626),
    .X(_0532_));
 sg13g2_a22oi_1 _3060_ (.Y(_0533_),
    .B1(_0532_),
    .B2(net589),
    .A2(_0444_),
    .A1(net591));
 sg13g2_nand4_1 _3061_ (.B(_0526_),
    .C(_0528_),
    .A(_0525_),
    .Y(_0534_),
    .D(_0533_));
 sg13g2_a221oi_1 _3062_ (.B2(net593),
    .C1(_0534_),
    .B1(_0523_),
    .A1(net598),
    .Y(_0535_),
    .A2(_0436_));
 sg13g2_or3_1 _3063_ (.A(net843),
    .B(_0514_),
    .C(_0535_),
    .X(_0536_));
 sg13g2_o21ai_1 _3064_ (.B1(_0536_),
    .Y(uio_out[3]),
    .A1(_0489_),
    .A2(_0490_));
 sg13g2_nand3_1 _3065_ (.B(_0462_),
    .C(_0463_),
    .A(net600),
    .Y(_0537_));
 sg13g2_nand3_1 _3066_ (.B(_0456_),
    .C(_0457_),
    .A(net804),
    .Y(_0538_));
 sg13g2_nand3_1 _3067_ (.B(_1510_),
    .C(_1511_),
    .A(net643),
    .Y(_0539_));
 sg13g2_nand3_1 _3068_ (.B(_0538_),
    .C(_0539_),
    .A(net637),
    .Y(_0540_));
 sg13g2_nand3_1 _3069_ (.B(_0458_),
    .C(_0459_),
    .A(net810),
    .Y(_0541_));
 sg13g2_nand3_1 _3070_ (.B(_0460_),
    .C(_0461_),
    .A(net819),
    .Y(_0542_));
 sg13g2_nand3_1 _3071_ (.B(_0540_),
    .C(_0541_),
    .A(net630),
    .Y(_0543_));
 sg13g2_nand3_1 _3072_ (.B(_0542_),
    .C(_0543_),
    .A(net595),
    .Y(_0544_));
 sg13g2_a21oi_1 _3073_ (.A1(_1132_),
    .A2(_1133_),
    .Y(_0545_),
    .B1(net602));
 sg13g2_a22oi_1 _3074_ (.Y(_0546_),
    .B1(net620),
    .B2(net762),
    .A2(net623),
    .A1(net716));
 sg13g2_a21oi_1 _3075_ (.A1(net726),
    .A2(net614),
    .Y(_0547_),
    .B1(net849));
 sg13g2_and2_1 _3076_ (.A(net841),
    .B(\a[21] ),
    .X(_0548_));
 sg13g2_nor2_1 _3077_ (.A(net834),
    .B(_0548_),
    .Y(_0549_));
 sg13g2_a21oi_1 _3078_ (.A1(\a[20] ),
    .A2(_0548_),
    .Y(_0550_),
    .B1(net835));
 sg13g2_o21ai_1 _3079_ (.B1(_0550_),
    .Y(_0551_),
    .A1(\a[20] ),
    .A2(\a[21] ));
 sg13g2_and2_1 _3080_ (.A(_1406_),
    .B(_0548_),
    .X(_0552_));
 sg13g2_o21ai_1 _3081_ (.B1(\a[20] ),
    .Y(_0553_),
    .A1(net610),
    .A2(_0552_));
 sg13g2_nand4_1 _3082_ (.B(_0547_),
    .C(_0551_),
    .A(_0546_),
    .Y(_0554_),
    .D(_0553_));
 sg13g2_nor2_1 _3083_ (.A(_0545_),
    .B(_0554_),
    .Y(_0555_));
 sg13g2_nand3_1 _3084_ (.B(_0544_),
    .C(_0555_),
    .A(_0537_),
    .Y(_0556_));
 sg13g2_or3_1 _3085_ (.A(_1153_),
    .B(_1154_),
    .C(net602),
    .X(_0557_));
 sg13g2_a22oi_1 _3086_ (.Y(_0558_),
    .B1(net837),
    .B2(_0482_),
    .A2(net605),
    .A1(\a[28] ));
 sg13g2_nor2b_1 _3087_ (.A(_0558_),
    .B_N(\a[29] ),
    .Y(_0559_));
 sg13g2_o21ai_1 _3088_ (.B1(net607),
    .Y(_0560_),
    .A1(\a[29] ),
    .A2(net836));
 sg13g2_a22oi_1 _3089_ (.Y(_0561_),
    .B1(net615),
    .B2(\ayayayayayaya.b[28] ),
    .A2(net624),
    .A1(\ayayayayayaya.b[30] ));
 sg13g2_a221oi_1 _3090_ (.B2(\a[28] ),
    .C1(_0559_),
    .B1(_0560_),
    .A1(net745),
    .Y(_0562_),
    .A2(net619));
 sg13g2_nand4_1 _3091_ (.B(_0557_),
    .C(_0561_),
    .A(net848),
    .Y(_0563_),
    .D(_0562_));
 sg13g2_nor3_1 _3092_ (.A(net650),
    .B(net645),
    .C(_0378_),
    .Y(_0564_));
 sg13g2_nor2_1 _3093_ (.A(net813),
    .B(_0564_),
    .Y(_0565_));
 sg13g2_a21oi_1 _3094_ (.A1(_0474_),
    .A2(_0475_),
    .Y(_0566_),
    .B1(net636));
 sg13g2_nor3_1 _3095_ (.A(net820),
    .B(_0565_),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_a21o_1 _3096_ (.A2(_0478_),
    .A1(net820),
    .B1(_0567_),
    .X(_0568_));
 sg13g2_a221oi_1 _3097_ (.B2(net596),
    .C1(_0563_),
    .B1(_0568_),
    .A1(net601),
    .Y(_0569_),
    .A2(_0479_));
 sg13g2_nor2_1 _3098_ (.A(_0600_),
    .B(_0569_),
    .Y(_0570_));
 sg13g2_nand3_1 _3099_ (.B(_0491_),
    .C(_0492_),
    .A(net804),
    .Y(_0571_));
 sg13g2_nand3_1 _3100_ (.B(_1361_),
    .C(_1362_),
    .A(net643),
    .Y(_0572_));
 sg13g2_nand3_1 _3101_ (.B(_0571_),
    .C(_0572_),
    .A(net638),
    .Y(_0573_));
 sg13g2_nand3_1 _3102_ (.B(_0493_),
    .C(_0494_),
    .A(net810),
    .Y(_0574_));
 sg13g2_a21oi_1 _3103_ (.A1(_0573_),
    .A2(_0574_),
    .Y(_0575_),
    .B1(net818));
 sg13g2_a21oi_1 _3104_ (.A1(_0495_),
    .A2(_0496_),
    .Y(_0576_),
    .B1(net630));
 sg13g2_or2_1 _3105_ (.X(_0577_),
    .B(_0576_),
    .A(_0575_));
 sg13g2_and3_2 _3106_ (.X(_0578_),
    .A(net794),
    .B(net801),
    .C(_0418_));
 sg13g2_mux2_1 _3107_ (.A0(_0509_),
    .A1(_0578_),
    .S(net635),
    .X(_0579_));
 sg13g2_mux2_1 _3108_ (.A0(_0510_),
    .A1(_0579_),
    .S(net629),
    .X(_0580_));
 sg13g2_o21ai_1 _3109_ (.B1(\a[13] ),
    .Y(_0581_),
    .A1(_0503_),
    .A2(_0505_));
 sg13g2_nor2_1 _3110_ (.A(\a[13] ),
    .B(net833),
    .Y(_0582_));
 sg13g2_o21ai_1 _3111_ (.B1(\a[12] ),
    .Y(_0583_),
    .A1(net609),
    .A2(_0582_));
 sg13g2_a22oi_1 _3112_ (.Y(_0584_),
    .B1(net619),
    .B2(net785),
    .A2(net625),
    .A1(net721));
 sg13g2_nand3_1 _3113_ (.B(_0581_),
    .C(_0583_),
    .A(net846),
    .Y(_0585_));
 sg13g2_a21oi_1 _3114_ (.A1(\ayayayayayaya.b[12] ),
    .A2(net612),
    .Y(_0586_),
    .B1(_0585_));
 sg13g2_a22oi_1 _3115_ (.Y(_0587_),
    .B1(_0580_),
    .B2(net590),
    .A2(_0511_),
    .A1(net592));
 sg13g2_nand3_1 _3116_ (.B(_0586_),
    .C(_0587_),
    .A(_0584_),
    .Y(_0588_));
 sg13g2_a221oi_1 _3117_ (.B2(net594),
    .C1(_0588_),
    .B1(_0577_),
    .A1(net599),
    .Y(_0589_),
    .A2(_0499_));
 sg13g2_nand3_1 _3118_ (.B(_0515_),
    .C(_0516_),
    .A(net800),
    .Y(_0590_));
 sg13g2_nand3_1 _3119_ (.B(_0103_),
    .C(_0104_),
    .A(net642),
    .Y(_0591_));
 sg13g2_nand3_1 _3120_ (.B(_0590_),
    .C(_0591_),
    .A(net633),
    .Y(_0592_));
 sg13g2_nand3_1 _3121_ (.B(_0517_),
    .C(_0518_),
    .A(net807),
    .Y(_0593_));
 sg13g2_a21oi_1 _3122_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0594_),
    .B1(net814));
 sg13g2_a21oi_1 _3123_ (.A1(_0519_),
    .A2(_0520_),
    .Y(_0595_),
    .B1(net626));
 sg13g2_or2_1 _3124_ (.X(_0596_),
    .B(_0595_),
    .A(_0594_));
 sg13g2_mux2_1 _3125_ (.A0(_0169_),
    .A1(_0529_),
    .S(net800),
    .X(_0597_));
 sg13g2_mux2_1 _3126_ (.A0(_0530_),
    .A1(_0597_),
    .S(net634),
    .X(_0598_));
 sg13g2_mux2_1 _3127_ (.A0(_0531_),
    .A1(_0598_),
    .S(net626),
    .X(_0599_));
 sg13g2_a21o_1 _3128_ (.A2(net623),
    .A1(net730),
    .B1(net849),
    .X(_0601_));
 sg13g2_a221oi_1 _3129_ (.B2(net795),
    .C1(_0601_),
    .B1(net611),
    .A1(net808),
    .Y(_0602_),
    .A2(net617));
 sg13g2_and2_1 _3130_ (.A(\a[5] ),
    .B(net604),
    .X(_0603_));
 sg13g2_o21ai_1 _3131_ (.B1(\a[4] ),
    .Y(_0604_),
    .A1(net608),
    .A2(_0603_));
 sg13g2_a21oi_1 _3132_ (.A1(net839),
    .A2(\a[5] ),
    .Y(_0605_),
    .B1(net832));
 sg13g2_or2_1 _3133_ (.X(_0606_),
    .B(\a[5] ),
    .A(\a[4] ));
 sg13g2_o21ai_1 _3134_ (.B1(_0606_),
    .Y(_0607_),
    .A1(_0527_),
    .A2(_0605_));
 sg13g2_a22oi_1 _3135_ (.Y(_0608_),
    .B1(_0599_),
    .B2(net589),
    .A2(_0532_),
    .A1(net591));
 sg13g2_nand4_1 _3136_ (.B(_0604_),
    .C(_0607_),
    .A(_0602_),
    .Y(_0609_),
    .D(_0608_));
 sg13g2_a221oi_1 _3137_ (.B2(net593),
    .C1(_0609_),
    .B1(_0596_),
    .A1(net598),
    .Y(_0610_),
    .A2(_0523_));
 sg13g2_nor3_1 _3138_ (.A(net843),
    .B(_0589_),
    .C(_0610_),
    .Y(_0612_));
 sg13g2_a21o_2 _3139_ (.A2(_0570_),
    .A1(_0556_),
    .B1(_0612_),
    .X(uio_out[4]));
 sg13g2_nand2_1 _3140_ (.Y(_0613_),
    .A(\a[30] ),
    .B(net625));
 sg13g2_a22oi_1 _3141_ (.Y(_0614_),
    .B1(net614),
    .B2(\ayayayayayaya.b[29] ),
    .A2(net619),
    .A1(\a[14] ));
 sg13g2_nand2_1 _3142_ (.Y(_0615_),
    .A(net841),
    .B(\a[30] ));
 sg13g2_o21ai_1 _3143_ (.B1(net607),
    .Y(_0616_),
    .A1(_1407_),
    .A2(_0615_));
 sg13g2_nand2_1 _3144_ (.Y(_0617_),
    .A(_1416_),
    .B(_0615_));
 sg13g2_o21ai_1 _3145_ (.B1(_0617_),
    .Y(_0618_),
    .A1(\a[29] ),
    .A2(net836));
 sg13g2_o21ai_1 _3146_ (.B1(_0618_),
    .Y(_0619_),
    .A1(\a[29] ),
    .A2(\a[30] ));
 sg13g2_nand4_1 _3147_ (.B(_0613_),
    .C(_0614_),
    .A(net849),
    .Y(_0620_),
    .D(_0619_));
 sg13g2_a221oi_1 _3148_ (.B2(\a[29] ),
    .C1(_0620_),
    .B1(_0616_),
    .A1(_1201_),
    .Y(_0622_),
    .A2(_1423_));
 sg13g2_a21o_1 _3149_ (.A2(_0564_),
    .A1(net813),
    .B1(net821),
    .X(_0623_));
 sg13g2_o21ai_1 _3150_ (.B1(net820),
    .Y(_0624_),
    .A1(_0565_),
    .A2(_0566_));
 sg13g2_nand3_1 _3151_ (.B(_0623_),
    .C(_0624_),
    .A(net596),
    .Y(_0625_));
 sg13g2_nand2_1 _3152_ (.Y(_0626_),
    .A(_0622_),
    .B(_0625_));
 sg13g2_a21oi_1 _3153_ (.A1(net601),
    .A2(_0568_),
    .Y(_0627_),
    .B1(_0626_));
 sg13g2_nand3_1 _3154_ (.B(_1512_),
    .C(_1517_),
    .A(net637),
    .Y(_0628_));
 sg13g2_nand3_1 _3155_ (.B(_0538_),
    .C(_0539_),
    .A(net810),
    .Y(_0629_));
 sg13g2_nand3_1 _3156_ (.B(_0540_),
    .C(_0541_),
    .A(net818),
    .Y(_0630_));
 sg13g2_nand3_1 _3157_ (.B(_0628_),
    .C(_0629_),
    .A(net630),
    .Y(_0631_));
 sg13g2_nand3_1 _3158_ (.B(_0630_),
    .C(_0631_),
    .A(net595),
    .Y(_0633_));
 sg13g2_nand3_1 _3159_ (.B(_0542_),
    .C(_0543_),
    .A(net600),
    .Y(_0634_));
 sg13g2_a21oi_1 _3160_ (.A1(\a[26] ),
    .A2(net624),
    .Y(_0635_),
    .B1(net848));
 sg13g2_a22oi_1 _3161_ (.Y(_0636_),
    .B1(net613),
    .B2(net724),
    .A2(net618),
    .A1(\a[10] ));
 sg13g2_o21ai_1 _3162_ (.B1(\a[22] ),
    .Y(_0637_),
    .A1(_0549_),
    .A2(_0552_));
 sg13g2_nor2_1 _3163_ (.A(\a[22] ),
    .B(net835),
    .Y(_0638_));
 sg13g2_o21ai_1 _3164_ (.B1(\a[21] ),
    .Y(_0639_),
    .A1(_1410_),
    .A2(_0638_));
 sg13g2_nand4_1 _3165_ (.B(_0636_),
    .C(_0637_),
    .A(_0635_),
    .Y(_0640_),
    .D(_0639_));
 sg13g2_a21oi_1 _3166_ (.A1(_1090_),
    .A2(_1091_),
    .Y(_0641_),
    .B1(net603));
 sg13g2_nor2_1 _3167_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sg13g2_nand3_1 _3168_ (.B(_0634_),
    .C(_0642_),
    .A(_0633_),
    .Y(_0644_));
 sg13g2_nand2_1 _3169_ (.Y(_0645_),
    .A(net844),
    .B(_0644_));
 sg13g2_nand3_1 _3170_ (.B(_1363_),
    .C(_1364_),
    .A(net638),
    .Y(_0646_));
 sg13g2_nand3_1 _3171_ (.B(_0571_),
    .C(_0572_),
    .A(net810),
    .Y(_0647_));
 sg13g2_a21oi_1 _3172_ (.A1(_0646_),
    .A2(_0647_),
    .Y(_0648_),
    .B1(net818));
 sg13g2_a21oi_1 _3173_ (.A1(_0573_),
    .A2(_0574_),
    .Y(_0649_),
    .B1(net630));
 sg13g2_or2_1 _3174_ (.X(_0650_),
    .B(_0649_),
    .A(_0648_));
 sg13g2_nand3_1 _3175_ (.B(net629),
    .C(_0578_),
    .A(net809),
    .Y(_0651_));
 sg13g2_nand2_1 _3176_ (.Y(_0652_),
    .A(net815),
    .B(_0579_));
 sg13g2_nand2_1 _3177_ (.Y(_0653_),
    .A(_0651_),
    .B(_0652_));
 sg13g2_and2_1 _3178_ (.A(\a[14] ),
    .B(net605),
    .X(_0655_));
 sg13g2_o21ai_1 _3179_ (.B1(\a[13] ),
    .Y(_0656_),
    .A1(net609),
    .A2(_0655_));
 sg13g2_a21oi_1 _3180_ (.A1(net840),
    .A2(\a[14] ),
    .Y(_0657_),
    .B1(net833));
 sg13g2_or2_1 _3181_ (.X(_0658_),
    .B(\a[14] ),
    .A(\a[13] ));
 sg13g2_o21ai_1 _3182_ (.B1(_0658_),
    .Y(_0659_),
    .A1(_0582_),
    .A2(_0657_));
 sg13g2_a22oi_1 _3183_ (.Y(_0660_),
    .B1(net616),
    .B2(\a[6] ),
    .A2(net621),
    .A1(\a[22] ));
 sg13g2_inv_1 _3184_ (.Y(_0661_),
    .A(_0660_));
 sg13g2_a221oi_1 _3185_ (.B2(_0653_),
    .C1(_0661_),
    .B1(net590),
    .A1(net748),
    .Y(_0662_),
    .A2(net612));
 sg13g2_nand4_1 _3186_ (.B(_0656_),
    .C(_0659_),
    .A(net846),
    .Y(_0663_),
    .D(_0662_));
 sg13g2_a21o_1 _3187_ (.A2(_0580_),
    .A1(net592),
    .B1(_0663_),
    .X(_0664_));
 sg13g2_a221oi_1 _3188_ (.B2(net594),
    .C1(_0664_),
    .B1(_0650_),
    .A1(net599),
    .Y(_0666_),
    .A2(_0577_));
 sg13g2_nand3_1 _3189_ (.B(_0105_),
    .C(_0106_),
    .A(net635),
    .Y(_0667_));
 sg13g2_nand3_1 _3190_ (.B(_0590_),
    .C(_0591_),
    .A(net807),
    .Y(_0668_));
 sg13g2_a21oi_1 _3191_ (.A1(_0667_),
    .A2(_0668_),
    .Y(_0669_),
    .B1(net814));
 sg13g2_a21oi_1 _3192_ (.A1(_0592_),
    .A2(_0593_),
    .Y(_0670_),
    .B1(net628));
 sg13g2_or2_1 _3193_ (.X(_0671_),
    .B(_0670_),
    .A(_0669_));
 sg13g2_a21o_1 _3194_ (.A2(net616),
    .A1(\a[2] ),
    .B1(net845),
    .X(_0672_));
 sg13g2_a221oi_1 _3195_ (.B2(net788),
    .C1(_0672_),
    .B1(net612),
    .A1(\a[18] ),
    .Y(_0673_),
    .A2(net621));
 sg13g2_o21ai_1 _3196_ (.B1(\a[6] ),
    .Y(_0674_),
    .A1(_0603_),
    .A2(_0605_));
 sg13g2_nor2_1 _3197_ (.A(\a[6] ),
    .B(net832),
    .Y(_0675_));
 sg13g2_o21ai_1 _3198_ (.B1(\a[5] ),
    .Y(_0677_),
    .A1(net608),
    .A2(_0675_));
 sg13g2_mux2_1 _3199_ (.A0(_0170_),
    .A1(_0597_),
    .S(net807),
    .X(_0678_));
 sg13g2_mux2_1 _3200_ (.A0(_0598_),
    .A1(_0678_),
    .S(net626),
    .X(_0679_));
 sg13g2_a22oi_1 _3201_ (.Y(_0680_),
    .B1(_0679_),
    .B2(net590),
    .A2(_0599_),
    .A1(net592));
 sg13g2_nand4_1 _3202_ (.B(_0674_),
    .C(_0677_),
    .A(_0673_),
    .Y(_0681_),
    .D(_0680_));
 sg13g2_a221oi_1 _3203_ (.B2(net593),
    .C1(_0681_),
    .B1(_0671_),
    .A1(net598),
    .Y(_0682_),
    .A2(_0596_));
 sg13g2_or3_1 _3204_ (.A(net843),
    .B(_0666_),
    .C(_0682_),
    .X(_0683_));
 sg13g2_o21ai_1 _3205_ (.B1(_0683_),
    .Y(uio_out[5]),
    .A1(_0627_),
    .A2(_0645_));
 sg13g2_a21oi_1 _3206_ (.A1(_1522_),
    .A2(_1523_),
    .Y(_0684_),
    .B1(net818));
 sg13g2_a21oi_1 _3207_ (.A1(_0628_),
    .A2(_0629_),
    .Y(_0685_),
    .B1(net630));
 sg13g2_o21ai_1 _3208_ (.B1(net595),
    .Y(_0687_),
    .A1(_0684_),
    .A2(_0685_));
 sg13g2_nand3_1 _3209_ (.B(_0630_),
    .C(_0631_),
    .A(net600),
    .Y(_0688_));
 sg13g2_a21oi_1 _3210_ (.A1(net841),
    .A2(\a[23] ),
    .Y(_0689_),
    .B1(net835));
 sg13g2_o21ai_1 _3211_ (.B1(\a[22] ),
    .Y(_0690_),
    .A1(net610),
    .A2(_0689_));
 sg13g2_a21oi_1 _3212_ (.A1(net754),
    .A2(net620),
    .Y(_0691_),
    .B1(net848));
 sg13g2_a22oi_1 _3213_ (.Y(_0692_),
    .B1(net615),
    .B2(net721),
    .A2(net623),
    .A1(\ayayayayayaya.b[27] ));
 sg13g2_nand3_1 _3214_ (.B(_0691_),
    .C(_0692_),
    .A(_0690_),
    .Y(_0693_));
 sg13g2_a21o_1 _3215_ (.A2(net605),
    .A1(\a[22] ),
    .B1(_0638_),
    .X(_0694_));
 sg13g2_a221oi_1 _3216_ (.B2(\a[23] ),
    .C1(_0693_),
    .B1(_0694_),
    .A1(_1054_),
    .Y(_0695_),
    .A2(_1423_));
 sg13g2_nand3_1 _3217_ (.B(_0688_),
    .C(_0695_),
    .A(_0687_),
    .Y(_0696_));
 sg13g2_nand3_1 _3218_ (.B(_0623_),
    .C(_0624_),
    .A(net601),
    .Y(_0698_));
 sg13g2_a22oi_1 _3219_ (.Y(_0699_),
    .B1(_1416_),
    .B2(_0615_),
    .A2(net605),
    .A1(\a[30] ));
 sg13g2_o21ai_1 _3220_ (.B1(net606),
    .Y(_0700_),
    .A1(net829),
    .A2(net836));
 sg13g2_and3_1 _3221_ (.X(_0701_),
    .A(net813),
    .B(net821),
    .C(_0564_));
 sg13g2_a22oi_1 _3222_ (.Y(_0702_),
    .B1(_0700_),
    .B2(\a[30] ),
    .A2(net619),
    .A1(net741));
 sg13g2_o21ai_1 _3223_ (.B1(_0702_),
    .Y(_0703_),
    .A1(_0665_),
    .A2(_0699_));
 sg13g2_a221oi_1 _3224_ (.B2(\ayayayayayaya.b[30] ),
    .C1(_0703_),
    .B1(net614),
    .A1(\ayayayayayaya.b[31] ),
    .Y(_0704_),
    .A2(net625));
 sg13g2_a22oi_1 _3225_ (.Y(_0705_),
    .B1(_0701_),
    .B2(net596),
    .A2(_1423_),
    .A1(_1253_));
 sg13g2_nand4_1 _3226_ (.B(_0698_),
    .C(_0704_),
    .A(net849),
    .Y(_0706_),
    .D(_0705_));
 sg13g2_nand3_1 _3227_ (.B(_0696_),
    .C(_0706_),
    .A(net844),
    .Y(_0707_));
 sg13g2_nand3_1 _3228_ (.B(_0667_),
    .C(_0668_),
    .A(net814),
    .Y(_0709_));
 sg13g2_nand3_1 _3229_ (.B(_0107_),
    .C(_0108_),
    .A(net629),
    .Y(_0710_));
 sg13g2_and2_1 _3230_ (.A(_0709_),
    .B(_0710_),
    .X(_0711_));
 sg13g2_a21oi_1 _3231_ (.A1(\a[6] ),
    .A2(net604),
    .Y(_0712_),
    .B1(_0675_));
 sg13g2_nand2b_1 _3232_ (.Y(_0713_),
    .B(net826),
    .A_N(_0712_));
 sg13g2_a21oi_1 _3233_ (.A1(net839),
    .A2(net826),
    .Y(_0714_),
    .B1(net832));
 sg13g2_o21ai_1 _3234_ (.B1(\a[6] ),
    .Y(_0715_),
    .A1(net608),
    .A2(_0714_));
 sg13g2_a22oi_1 _3235_ (.Y(_0716_),
    .B1(net611),
    .B2(net785),
    .A2(net621),
    .A1(\ayayayayayaya.b[19] ));
 sg13g2_a21oi_1 _3236_ (.A1(\ayayayayayaya.b[3] ),
    .A2(net616),
    .Y(_0717_),
    .B1(net845));
 sg13g2_nand4_1 _3237_ (.B(_0715_),
    .C(_0716_),
    .A(_0713_),
    .Y(_0718_),
    .D(_0717_));
 sg13g2_mux2_1 _3238_ (.A0(_0171_),
    .A1(_0678_),
    .S(net814),
    .X(_0720_));
 sg13g2_a221oi_1 _3239_ (.B2(net591),
    .C1(_0718_),
    .B1(_0679_),
    .A1(net598),
    .Y(_0721_),
    .A2(_0671_));
 sg13g2_a22oi_1 _3240_ (.Y(_0722_),
    .B1(_0720_),
    .B2(net589),
    .A2(_0711_),
    .A1(net593));
 sg13g2_nand3_1 _3241_ (.B(_0646_),
    .C(_0647_),
    .A(net818),
    .Y(_0723_));
 sg13g2_nand3_1 _3242_ (.B(_1365_),
    .C(_1366_),
    .A(net630),
    .Y(_0724_));
 sg13g2_nand3_1 _3243_ (.B(_0723_),
    .C(_0724_),
    .A(net596),
    .Y(_0725_));
 sg13g2_nand2_1 _3244_ (.Y(_0726_),
    .A(net592),
    .B(_0653_));
 sg13g2_nand2_1 _3245_ (.Y(_0727_),
    .A(net745),
    .B(net612));
 sg13g2_o21ai_1 _3246_ (.B1(net824),
    .Y(_0728_),
    .A1(_0655_),
    .A2(_0657_));
 sg13g2_nor2_1 _3247_ (.A(net824),
    .B(_1417_),
    .Y(_0729_));
 sg13g2_o21ai_1 _3248_ (.B1(\a[14] ),
    .Y(_0731_),
    .A1(net609),
    .A2(_0729_));
 sg13g2_nand4_1 _3249_ (.B(_0727_),
    .C(_0728_),
    .A(net846),
    .Y(_0732_),
    .D(_0731_));
 sg13g2_a221oi_1 _3250_ (.B2(net779),
    .C1(_0732_),
    .B1(net618),
    .A1(net720),
    .Y(_0733_),
    .A2(net622));
 sg13g2_nand4_1 _3251_ (.B(net817),
    .C(net590),
    .A(net808),
    .Y(_0734_),
    .D(_0578_));
 sg13g2_nand4_1 _3252_ (.B(_0726_),
    .C(_0733_),
    .A(_0725_),
    .Y(_0735_),
    .D(_0734_));
 sg13g2_a21oi_1 _3253_ (.A1(net598),
    .A2(_0650_),
    .Y(_0736_),
    .B1(_0735_));
 sg13g2_a21o_1 _3254_ (.A2(_0722_),
    .A1(_0721_),
    .B1(net843),
    .X(_0737_));
 sg13g2_o21ai_1 _3255_ (.B1(_0707_),
    .Y(uio_out[6]),
    .A1(_0736_),
    .A2(_0737_));
 sg13g2_nand3_1 _3256_ (.B(_1368_),
    .C(net595),
    .A(_1367_),
    .Y(_0738_));
 sg13g2_nand3_1 _3257_ (.B(_0723_),
    .C(_0724_),
    .A(net601),
    .Y(_0739_));
 sg13g2_nand4_1 _3258_ (.B(net814),
    .C(net592),
    .A(net809),
    .Y(_0741_),
    .D(_0578_));
 sg13g2_nand3_1 _3259_ (.B(net830),
    .C(net604),
    .A(net1),
    .Y(_0742_));
 sg13g2_nand3_1 _3260_ (.B(net838),
    .C(_1422_),
    .A(net827),
    .Y(_0743_));
 sg13g2_nand3_1 _3261_ (.B(_0742_),
    .C(_0743_),
    .A(net606),
    .Y(_0744_));
 sg13g2_nand2_1 _3262_ (.Y(_0745_),
    .A(_1401_),
    .B(net837));
 sg13g2_nand3_1 _3263_ (.B(net1),
    .C(net837),
    .A(net840),
    .Y(_0746_));
 sg13g2_and2_1 _3264_ (.A(net824),
    .B(net830),
    .X(_0747_));
 sg13g2_o21ai_1 _3265_ (.B1(_0745_),
    .Y(_0748_),
    .A1(_0746_),
    .A2(_0747_));
 sg13g2_o21ai_1 _3266_ (.B1(_0748_),
    .Y(_0749_),
    .A1(net824),
    .A2(net830));
 sg13g2_nand2_1 _3267_ (.Y(_0750_),
    .A(net826),
    .B(net617));
 sg13g2_a22oi_1 _3268_ (.Y(_0752_),
    .B1(net613),
    .B2(net741),
    .A2(net622),
    .A1(\a[23] ));
 sg13g2_or2_1 _3269_ (.X(_0753_),
    .B(net824),
    .A(net827));
 sg13g2_nand2_1 _3270_ (.Y(_0754_),
    .A(_1403_),
    .B(net837));
 sg13g2_nand2_1 _3271_ (.Y(_0755_),
    .A(net837),
    .B(_1422_));
 sg13g2_and2_1 _3272_ (.A(net827),
    .B(\a[15] ),
    .X(_0756_));
 sg13g2_o21ai_1 _3273_ (.B1(_0754_),
    .Y(_0757_),
    .A1(_0755_),
    .A2(_0756_));
 sg13g2_nand4_1 _3274_ (.B(_0749_),
    .C(_0750_),
    .A(net846),
    .Y(_0758_),
    .D(_0752_));
 sg13g2_a221oi_1 _3275_ (.B2(_0757_),
    .C1(_0758_),
    .B1(_0753_),
    .A1(\a[15] ),
    .Y(_0759_),
    .A2(_0744_));
 sg13g2_nand4_1 _3276_ (.B(_0739_),
    .C(_0741_),
    .A(_0738_),
    .Y(_0760_),
    .D(_0759_));
 sg13g2_nand3_1 _3277_ (.B(_0709_),
    .C(_0710_),
    .A(net598),
    .Y(_0761_));
 sg13g2_nand3_1 _3278_ (.B(_0109_),
    .C(_0110_),
    .A(net593),
    .Y(_0763_));
 sg13g2_nand2_1 _3279_ (.Y(_0764_),
    .A(net779),
    .B(net612));
 sg13g2_a22oi_1 _3280_ (.Y(_0765_),
    .B1(net617),
    .B2(\a[3] ),
    .A2(net621),
    .A1(\a[19] ));
 sg13g2_o21ai_1 _3281_ (.B1(net826),
    .Y(_0766_),
    .A1(net608),
    .A2(_0182_));
 sg13g2_nand3_1 _3282_ (.B(net826),
    .C(net825),
    .A(net839),
    .Y(_0767_));
 sg13g2_nor2_1 _3283_ (.A(net826),
    .B(net825),
    .Y(_0768_));
 sg13g2_nor2_1 _3284_ (.A(net833),
    .B(_0768_),
    .Y(_0769_));
 sg13g2_a21oi_1 _3285_ (.A1(_0767_),
    .A2(_0769_),
    .Y(_0770_),
    .B1(net847));
 sg13g2_nand4_1 _3286_ (.B(_0765_),
    .C(_0766_),
    .A(_0764_),
    .Y(_0771_),
    .D(_0770_));
 sg13g2_a221oi_1 _3287_ (.B2(net591),
    .C1(_0771_),
    .B1(_0720_),
    .A1(_0179_),
    .Y(_0772_),
    .A2(net589));
 sg13g2_nand3_1 _3288_ (.B(_0763_),
    .C(_0772_),
    .A(_0761_),
    .Y(_0774_));
 sg13g2_nand3_1 _3289_ (.B(_0760_),
    .C(_0774_),
    .A(_0600_),
    .Y(_0775_));
 sg13g2_nand3_1 _3290_ (.B(_1524_),
    .C(_1536_),
    .A(net595),
    .Y(_0776_));
 sg13g2_o21ai_1 _3291_ (.B1(net600),
    .Y(_0777_),
    .A1(_0684_),
    .A2(_0685_));
 sg13g2_nand3_1 _3292_ (.B(\a[23] ),
    .C(\a[24] ),
    .A(net841),
    .Y(_0778_));
 sg13g2_o21ai_1 _3293_ (.B1(_0778_),
    .Y(_0779_),
    .A1(\a[23] ),
    .A2(\a[24] ));
 sg13g2_nor2_1 _3294_ (.A(net836),
    .B(_0779_),
    .Y(_0780_));
 sg13g2_a21oi_1 _3295_ (.A1(\a[27] ),
    .A2(net625),
    .Y(_0781_),
    .B1(net848));
 sg13g2_a22oi_1 _3296_ (.Y(_0782_),
    .B1(net610),
    .B2(\a[23] ),
    .A2(net614),
    .A1(net720));
 sg13g2_nor2_1 _3297_ (.A(_1407_),
    .B(_0778_),
    .Y(_0783_));
 sg13g2_a21oi_1 _3298_ (.A1(\a[11] ),
    .A2(net618),
    .Y(_0785_),
    .B1(_0783_));
 sg13g2_nand3_1 _3299_ (.B(_0782_),
    .C(_0785_),
    .A(_0781_),
    .Y(_0786_));
 sg13g2_a21oi_1 _3300_ (.A1(_1019_),
    .A2(_1020_),
    .Y(_0787_),
    .B1(net602));
 sg13g2_nor3_1 _3301_ (.A(_0780_),
    .B(_0786_),
    .C(_0787_),
    .Y(_0788_));
 sg13g2_nand3_1 _3302_ (.B(_0777_),
    .C(_0788_),
    .A(_0776_),
    .Y(_0789_));
 sg13g2_nand3_1 _3303_ (.B(net838),
    .C(_1422_),
    .A(net831),
    .Y(_0790_));
 sg13g2_nand3_1 _3304_ (.B(net828),
    .C(net604),
    .A(net1),
    .Y(_0791_));
 sg13g2_nor2_1 _3305_ (.A(net622),
    .B(net609),
    .Y(_0792_));
 sg13g2_nand3_1 _3306_ (.B(_0791_),
    .C(_0792_),
    .A(_0790_),
    .Y(_0793_));
 sg13g2_and2_1 _3307_ (.A(net828),
    .B(net829),
    .X(_0794_));
 sg13g2_o21ai_1 _3308_ (.B1(_0745_),
    .Y(_0796_),
    .A1(_0746_),
    .A2(_0794_));
 sg13g2_o21ai_1 _3309_ (.B1(_0796_),
    .Y(_0797_),
    .A1(net827),
    .A2(net829));
 sg13g2_and2_1 _3310_ (.A(net830),
    .B(net829),
    .X(_0798_));
 sg13g2_o21ai_1 _3311_ (.B1(_0754_),
    .Y(_0799_),
    .A1(_0755_),
    .A2(_0798_));
 sg13g2_o21ai_1 _3312_ (.B1(_0799_),
    .Y(_0800_),
    .A1(net830),
    .A2(net829));
 sg13g2_a22oi_1 _3313_ (.Y(_0801_),
    .B1(net613),
    .B2(\ayayayayayaya.b[31] ),
    .A2(net618),
    .A1(net824));
 sg13g2_nand4_1 _3314_ (.B(_0797_),
    .C(_0800_),
    .A(net846),
    .Y(_0802_),
    .D(_0801_));
 sg13g2_a21oi_1 _3315_ (.A1(net829),
    .A2(_0793_),
    .Y(_0803_),
    .B1(_0802_));
 sg13g2_a22oi_1 _3316_ (.Y(_0804_),
    .B1(_0701_),
    .B2(net601),
    .A2(_1423_),
    .A1(_1308_));
 sg13g2_a21oi_1 _3317_ (.A1(_0803_),
    .A2(_0804_),
    .Y(_0805_),
    .B1(_0600_));
 sg13g2_nand2_1 _3318_ (.Y(_0807_),
    .A(_0789_),
    .B(_0805_));
 sg13g2_nand2_2 _3319_ (.Y(uio_out[7]),
    .A(_0775_),
    .B(_0807_));
 sg13g2_nand2b_1 _3320_ (.Y(_0808_),
    .B(net844),
    .A_N(net846));
 sg13g2_nor3_2 _3321_ (.A(net5),
    .B(net606),
    .C(_0808_),
    .Y(_0809_));
 sg13g2_mux2_1 _3322_ (.A0(net830),
    .A1(net6),
    .S(_0809_),
    .X(_0000_));
 sg13g2_mux2_1 _3323_ (.A0(net107),
    .A1(net7),
    .S(_0809_),
    .X(_0001_));
 sg13g2_mux2_1 _3324_ (.A0(net112),
    .A1(net8),
    .S(_0809_),
    .X(_0002_));
 sg13g2_mux2_1 _3325_ (.A0(net97),
    .A1(net9),
    .S(_0809_),
    .X(_0003_));
 sg13g2_mux2_1 _3326_ (.A0(net110),
    .A1(net10),
    .S(_0809_),
    .X(_0004_));
 sg13g2_mux2_1 _3327_ (.A0(net98),
    .A1(net11),
    .S(_0809_),
    .X(_0005_));
 sg13g2_mux2_1 _3328_ (.A0(net109),
    .A1(net12),
    .S(_0809_),
    .X(_0006_));
 sg13g2_mux2_1 _3329_ (.A0(net106),
    .A1(net13),
    .S(_0809_),
    .X(_0007_));
 sg13g2_nand2_1 _3330_ (.Y(_0811_),
    .A(net844),
    .B(net846));
 sg13g2_nor3_2 _3331_ (.A(net5),
    .B(net606),
    .C(_0811_),
    .Y(_0812_));
 sg13g2_mux2_1 _3332_ (.A0(net92),
    .A1(net6),
    .S(net588),
    .X(_0008_));
 sg13g2_mux2_1 _3333_ (.A0(net90),
    .A1(net7),
    .S(net588),
    .X(_0009_));
 sg13g2_mux2_1 _3334_ (.A0(net84),
    .A1(net8),
    .S(net588),
    .X(_0010_));
 sg13g2_mux2_1 _3335_ (.A0(net89),
    .A1(net9),
    .S(net588),
    .X(_0011_));
 sg13g2_mux2_1 _3336_ (.A0(net102),
    .A1(net10),
    .S(_0812_),
    .X(_0012_));
 sg13g2_mux2_1 _3337_ (.A0(net96),
    .A1(net11),
    .S(net588),
    .X(_0013_));
 sg13g2_mux2_1 _3338_ (.A0(net88),
    .A1(net12),
    .S(net588),
    .X(_0014_));
 sg13g2_nand2_1 _3339_ (.Y(_0814_),
    .A(net13),
    .B(net588));
 sg13g2_o21ai_1 _3340_ (.B1(_0814_),
    .Y(_0015_),
    .A1(_0665_),
    .A2(net588));
 sg13g2_nor4_2 _3341_ (.A(net5),
    .B(net844),
    .C(net847),
    .Y(_0815_),
    .D(net606));
 sg13g2_mux2_1 _3342_ (.A0(net78),
    .A1(net6),
    .S(net587),
    .X(_0016_));
 sg13g2_nand2_1 _3343_ (.Y(_0816_),
    .A(net7),
    .B(net587));
 sg13g2_o21ai_1 _3344_ (.B1(_0816_),
    .Y(_0017_),
    .A1(_0621_),
    .A2(net587));
 sg13g2_mux2_1 _3345_ (.A0(net95),
    .A1(net8),
    .S(_0815_),
    .X(_0018_));
 sg13g2_nand2_1 _3346_ (.Y(_0817_),
    .A(net9),
    .B(net587));
 sg13g2_o21ai_1 _3347_ (.B1(_0817_),
    .Y(_0019_),
    .A1(_0632_),
    .A2(net587));
 sg13g2_mux2_1 _3348_ (.A0(net105),
    .A1(net10),
    .S(_0815_),
    .X(_0020_));
 sg13g2_nand2_1 _3349_ (.Y(_0819_),
    .A(net11),
    .B(net587));
 sg13g2_o21ai_1 _3350_ (.B1(_0819_),
    .Y(_0021_),
    .A1(_0643_),
    .A2(net587));
 sg13g2_mux2_1 _3351_ (.A0(net103),
    .A1(net12),
    .S(net587),
    .X(_0022_));
 sg13g2_mux2_1 _3352_ (.A0(net79),
    .A1(net13),
    .S(_0815_),
    .X(_0023_));
 sg13g2_nand2_2 _3353_ (.Y(_0820_),
    .A(_0600_),
    .B(net845));
 sg13g2_nor3_2 _3354_ (.A(net5),
    .B(net606),
    .C(_0820_),
    .Y(_0821_));
 sg13g2_mux2_1 _3355_ (.A0(net80),
    .A1(net6),
    .S(net586),
    .X(_0024_));
 sg13g2_nand2_1 _3356_ (.Y(_0822_),
    .A(net7),
    .B(net586));
 sg13g2_o21ai_1 _3357_ (.B1(_0822_),
    .Y(_0025_),
    .A1(_0654_),
    .A2(net586));
 sg13g2_mux2_1 _3358_ (.A0(net93),
    .A1(net8),
    .S(net586),
    .X(_0026_));
 sg13g2_mux2_1 _3359_ (.A0(net94),
    .A1(net9),
    .S(net586),
    .X(_0027_));
 sg13g2_mux2_1 _3360_ (.A0(net108),
    .A1(net10),
    .S(net586),
    .X(_0028_));
 sg13g2_mux2_1 _3361_ (.A0(net104),
    .A1(net11),
    .S(net586),
    .X(_0029_));
 sg13g2_mux2_1 _3362_ (.A0(net99),
    .A1(net12),
    .S(_0821_),
    .X(_0030_));
 sg13g2_mux2_1 _3363_ (.A0(net83),
    .A1(net13),
    .S(net586),
    .X(_0031_));
 sg13g2_nor4_1 _3364_ (.A(net5),
    .B(net844),
    .C(net847),
    .D(_1409_),
    .Y(_0824_));
 sg13g2_mux2_1 _3365_ (.A0(net823),
    .A1(net6),
    .S(net585),
    .X(_0032_));
 sg13g2_nand2_1 _3366_ (.Y(_0825_),
    .A(net7),
    .B(net585));
 sg13g2_o21ai_1 _3367_ (.B1(_0825_),
    .Y(_0033_),
    .A1(net626),
    .A2(net585));
 sg13g2_nand2_1 _3368_ (.Y(_0827_),
    .A(net8),
    .B(net584));
 sg13g2_o21ai_1 _3369_ (.B1(_0827_),
    .Y(_0034_),
    .A1(net633),
    .A2(net585));
 sg13g2_nand2_1 _3370_ (.Y(_0828_),
    .A(net9),
    .B(net584));
 sg13g2_o21ai_1 _3371_ (.B1(_0828_),
    .Y(_0035_),
    .A1(net640),
    .A2(net585));
 sg13g2_nand2_1 _3372_ (.Y(_0829_),
    .A(net10),
    .B(net585));
 sg13g2_o21ai_1 _3373_ (.B1(_0829_),
    .Y(_0036_),
    .A1(net647),
    .A2(net585));
 sg13g2_nand2_1 _3374_ (.Y(_0830_),
    .A(net11),
    .B(net584));
 sg13g2_o21ai_1 _3375_ (.B1(_0830_),
    .Y(_0037_),
    .A1(net654),
    .A2(net584));
 sg13g2_nand2_1 _3376_ (.Y(_0831_),
    .A(net12),
    .B(net584));
 sg13g2_o21ai_1 _3377_ (.B1(_0831_),
    .Y(_0038_),
    .A1(net660),
    .A2(net584));
 sg13g2_nand2_1 _3378_ (.Y(_0833_),
    .A(net13),
    .B(net584));
 sg13g2_o21ai_1 _3379_ (.B1(_0833_),
    .Y(_0039_),
    .A1(net664),
    .A2(net584));
 sg13g2_nor3_2 _3380_ (.A(net5),
    .B(_1409_),
    .C(_0820_),
    .Y(_0834_));
 sg13g2_nand2_1 _3381_ (.Y(_0835_),
    .A(net6),
    .B(net582));
 sg13g2_o21ai_1 _3382_ (.B1(_0835_),
    .Y(_0040_),
    .A1(net670),
    .A2(net582));
 sg13g2_nand2_1 _3383_ (.Y(_0836_),
    .A(net7),
    .B(net582));
 sg13g2_o21ai_1 _3384_ (.B1(_0836_),
    .Y(_0041_),
    .A1(net676),
    .A2(net582));
 sg13g2_nand2_1 _3385_ (.Y(_0837_),
    .A(net8),
    .B(net582));
 sg13g2_o21ai_1 _3386_ (.B1(_0837_),
    .Y(_0042_),
    .A1(net679),
    .A2(net582));
 sg13g2_nand2_1 _3387_ (.Y(_0838_),
    .A(net9),
    .B(net582));
 sg13g2_o21ai_1 _3388_ (.B1(_0838_),
    .Y(_0043_),
    .A1(net682),
    .A2(net582));
 sg13g2_nand2_1 _3389_ (.Y(_0840_),
    .A(net10),
    .B(net583));
 sg13g2_o21ai_1 _3390_ (.B1(_0840_),
    .Y(_0044_),
    .A1(net686),
    .A2(net583));
 sg13g2_nand2_1 _3391_ (.Y(_0841_),
    .A(net11),
    .B(net583));
 sg13g2_o21ai_1 _3392_ (.B1(_0841_),
    .Y(_0045_),
    .A1(net689),
    .A2(net583));
 sg13g2_nand2_1 _3393_ (.Y(_0842_),
    .A(net12),
    .B(net583));
 sg13g2_o21ai_1 _3394_ (.B1(_0842_),
    .Y(_0046_),
    .A1(net693),
    .A2(net583));
 sg13g2_nand2_1 _3395_ (.Y(_0843_),
    .A(net13),
    .B(net583));
 sg13g2_o21ai_1 _3396_ (.B1(_0843_),
    .Y(_0047_),
    .A1(net697),
    .A2(net583));
 sg13g2_nor3_2 _3397_ (.A(net5),
    .B(_1409_),
    .C(_0808_),
    .Y(_0844_));
 sg13g2_nand2_1 _3398_ (.Y(_0846_),
    .A(net6),
    .B(net580));
 sg13g2_o21ai_1 _3399_ (.B1(_0846_),
    .Y(_0048_),
    .A1(net699),
    .A2(net580));
 sg13g2_nand2_1 _3400_ (.Y(_0847_),
    .A(net7),
    .B(net580));
 sg13g2_o21ai_1 _3401_ (.B1(_0847_),
    .Y(_0049_),
    .A1(net702),
    .A2(net580));
 sg13g2_nand2_1 _3402_ (.Y(_0848_),
    .A(net8),
    .B(net580));
 sg13g2_o21ai_1 _3403_ (.B1(_0848_),
    .Y(_0050_),
    .A1(net704),
    .A2(net580));
 sg13g2_nand2_1 _3404_ (.Y(_0849_),
    .A(net9),
    .B(net580));
 sg13g2_o21ai_1 _3405_ (.B1(_0849_),
    .Y(_0051_),
    .A1(net706),
    .A2(net580));
 sg13g2_nand2_1 _3406_ (.Y(_0850_),
    .A(net10),
    .B(net581));
 sg13g2_o21ai_1 _3407_ (.B1(_0850_),
    .Y(_0052_),
    .A1(net708),
    .A2(net581));
 sg13g2_nand2_1 _3408_ (.Y(_0852_),
    .A(net11),
    .B(net581));
 sg13g2_o21ai_1 _3409_ (.B1(_0852_),
    .Y(_0053_),
    .A1(net710),
    .A2(net581));
 sg13g2_nand2_1 _3410_ (.Y(_0853_),
    .A(net12),
    .B(net581));
 sg13g2_o21ai_1 _3411_ (.B1(_0853_),
    .Y(_0054_),
    .A1(net711),
    .A2(net581));
 sg13g2_nand2_1 _3412_ (.Y(_0854_),
    .A(net13),
    .B(net581));
 sg13g2_o21ai_1 _3413_ (.B1(_0854_),
    .Y(_0055_),
    .A1(_0740_),
    .A2(net581));
 sg13g2_nor3_1 _3414_ (.A(net5),
    .B(_1409_),
    .C(_0811_),
    .Y(_0855_));
 sg13g2_nand2_1 _3415_ (.Y(_0856_),
    .A(net6),
    .B(net579));
 sg13g2_o21ai_1 _3416_ (.B1(_0856_),
    .Y(_0056_),
    .A1(net714),
    .A2(net578));
 sg13g2_nand2_1 _3417_ (.Y(_0857_),
    .A(net7),
    .B(net579));
 sg13g2_o21ai_1 _3418_ (.B1(_0857_),
    .Y(_0057_),
    .A1(net715),
    .A2(net578));
 sg13g2_nand2_1 _3419_ (.Y(_0859_),
    .A(net8),
    .B(net579));
 sg13g2_o21ai_1 _3420_ (.B1(_0859_),
    .Y(_0058_),
    .A1(_0708_),
    .A2(net579));
 sg13g2_nand2_1 _3421_ (.Y(_0860_),
    .A(net9),
    .B(net579));
 sg13g2_o21ai_1 _3422_ (.B1(_0860_),
    .Y(_0059_),
    .A1(_0697_),
    .A2(net579));
 sg13g2_nand2_1 _3423_ (.Y(_0861_),
    .A(net10),
    .B(net578));
 sg13g2_o21ai_1 _3424_ (.B1(_0861_),
    .Y(_0060_),
    .A1(_0686_),
    .A2(net578));
 sg13g2_nand2_1 _3425_ (.Y(_0862_),
    .A(net11),
    .B(net578));
 sg13g2_o21ai_1 _3426_ (.B1(_0862_),
    .Y(_0061_),
    .A1(_0676_),
    .A2(net578));
 sg13g2_mux2_1 _3427_ (.A0(net85),
    .A1(net12),
    .S(net578),
    .X(_0062_));
 sg13g2_mux2_1 _3428_ (.A0(net86),
    .A1(net13),
    .S(net578),
    .X(_0063_));
 sg13g2_dfrbpq_1 _3429_ (.RESET_B(net68),
    .D(_0000_),
    .Q(\a[16] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _3430_ (.RESET_B(net67),
    .D(_0001_),
    .Q(\a[17] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _3431_ (.RESET_B(net66),
    .D(_0002_),
    .Q(\a[18] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _3432_ (.RESET_B(net65),
    .D(_0003_),
    .Q(\a[19] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _3433_ (.RESET_B(net64),
    .D(_0004_),
    .Q(\a[20] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _3434_ (.RESET_B(net63),
    .D(_0005_),
    .Q(\a[21] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _3435_ (.RESET_B(net62),
    .D(_0006_),
    .Q(\a[22] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _3436_ (.RESET_B(net61),
    .D(_0007_),
    .Q(\a[23] ),
    .CLK(clknet_4_6_0_clk));
 sg13g2_dfrbpq_2 _3437_ (.RESET_B(net60),
    .D(_0008_),
    .Q(\a[24] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _3438_ (.RESET_B(net59),
    .D(_0009_),
    .Q(\a[25] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _3439_ (.RESET_B(net58),
    .D(_0010_),
    .Q(\a[26] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _3440_ (.RESET_B(net57),
    .D(_0011_),
    .Q(\a[27] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _3441_ (.RESET_B(net56),
    .D(_0012_),
    .Q(\a[28] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _3442_ (.RESET_B(net55),
    .D(_0013_),
    .Q(\a[29] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _3443_ (.RESET_B(net54),
    .D(_0014_),
    .Q(\a[30] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _3444_ (.RESET_B(net53),
    .D(_0015_),
    .Q(\a[31] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_1 _3445_ (.RESET_B(net52),
    .D(_0016_),
    .Q(\a[0] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _3446_ (.RESET_B(net51),
    .D(_0017_),
    .Q(\a[1] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _3447_ (.RESET_B(net50),
    .D(_0018_),
    .Q(\a[2] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _3448_ (.RESET_B(net49),
    .D(_0019_),
    .Q(\a[3] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _3449_ (.RESET_B(net48),
    .D(_0020_),
    .Q(\a[4] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _3450_ (.RESET_B(net47),
    .D(_0021_),
    .Q(\a[5] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_2 _3451_ (.RESET_B(net46),
    .D(_0022_),
    .Q(\a[6] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _3452_ (.RESET_B(net45),
    .D(_0023_),
    .Q(\a[7] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_1 _3453_ (.RESET_B(net44),
    .D(_0024_),
    .Q(\a[8] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _3454_ (.RESET_B(net43),
    .D(_0025_),
    .Q(\a[9] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _3455_ (.RESET_B(net42),
    .D(_0026_),
    .Q(\a[10] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _3456_ (.RESET_B(net41),
    .D(_0027_),
    .Q(\a[11] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_2 _3457_ (.RESET_B(net40),
    .D(_0028_),
    .Q(\a[12] ),
    .CLK(clknet_4_7_0_clk));
 sg13g2_dfrbpq_2 _3458_ (.RESET_B(net39),
    .D(_0029_),
    .Q(\a[13] ),
    .CLK(clknet_4_4_0_clk));
 sg13g2_dfrbpq_2 _3459_ (.RESET_B(net38),
    .D(_0030_),
    .Q(\a[14] ),
    .CLK(clknet_4_3_0_clk));
 sg13g2_dfrbpq_2 _3460_ (.RESET_B(net37),
    .D(_0031_),
    .Q(\a[15] ),
    .CLK(clknet_4_5_0_clk));
 sg13g2_dfrbpq_1 _3461_ (.RESET_B(net36),
    .D(_0032_),
    .Q(\ayayayayayaya.b[0] ),
    .CLK(clknet_4_2_0_clk));
 sg13g2_dfrbpq_1 _3462_ (.RESET_B(net35),
    .D(_0033_),
    .Q(\ayayayayayaya.b[1] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_2 _3463_ (.RESET_B(net34),
    .D(_0034_),
    .Q(\ayayayayayaya.b[2] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_2 _3464_ (.RESET_B(net33),
    .D(_0035_),
    .Q(\ayayayayayaya.b[3] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _3465_ (.RESET_B(net32),
    .D(_0036_),
    .Q(\ayayayayayaya.b[4] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _3466_ (.RESET_B(net31),
    .D(_0037_),
    .Q(\ayayayayayaya.b[5] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _3467_ (.RESET_B(net30),
    .D(_0038_),
    .Q(\ayayayayayaya.b[6] ),
    .CLK(clknet_4_1_0_clk));
 sg13g2_dfrbpq_1 _3468_ (.RESET_B(net29),
    .D(_0039_),
    .Q(\ayayayayayaya.b[7] ),
    .CLK(clknet_4_0_0_clk));
 sg13g2_dfrbpq_1 _3469_ (.RESET_B(net28),
    .D(_0040_),
    .Q(\ayayayayayaya.b[8] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _3470_ (.RESET_B(net27),
    .D(_0041_),
    .Q(\ayayayayayaya.b[9] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_1 _3471_ (.RESET_B(net26),
    .D(_0042_),
    .Q(\ayayayayayaya.b[10] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _3472_ (.RESET_B(net25),
    .D(_0043_),
    .Q(\ayayayayayaya.b[11] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _3473_ (.RESET_B(net24),
    .D(_0044_),
    .Q(\ayayayayayaya.b[12] ),
    .CLK(clknet_4_11_0_clk));
 sg13g2_dfrbpq_2 _3474_ (.RESET_B(net23),
    .D(_0045_),
    .Q(\ayayayayayaya.b[13] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_2 _3475_ (.RESET_B(net22),
    .D(_0046_),
    .Q(\ayayayayayaya.b[14] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _3476_ (.RESET_B(net21),
    .D(_0047_),
    .Q(\ayayayayayaya.b[15] ),
    .CLK(clknet_4_10_0_clk));
 sg13g2_dfrbpq_1 _3477_ (.RESET_B(net20),
    .D(_0048_),
    .Q(\ayayayayayaya.b[16] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _3478_ (.RESET_B(net19),
    .D(_0049_),
    .Q(\ayayayayayaya.b[17] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _3479_ (.RESET_B(net18),
    .D(_0050_),
    .Q(\ayayayayayaya.b[18] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_2 _3480_ (.RESET_B(net17),
    .D(_0051_),
    .Q(\ayayayayayaya.b[19] ),
    .CLK(clknet_4_8_0_clk));
 sg13g2_dfrbpq_1 _3481_ (.RESET_B(net16),
    .D(_0052_),
    .Q(\ayayayayayaya.b[20] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _3482_ (.RESET_B(net15),
    .D(_0053_),
    .Q(\ayayayayayaya.b[21] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _3483_ (.RESET_B(net14),
    .D(_0054_),
    .Q(\ayayayayayaya.b[22] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_1 _3484_ (.RESET_B(net77),
    .D(_0055_),
    .Q(\ayayayayayaya.b[23] ),
    .CLK(clknet_4_15_0_clk));
 sg13g2_dfrbpq_2 _3485_ (.RESET_B(net76),
    .D(_0056_),
    .Q(\ayayayayayaya.b[24] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_1 _3486_ (.RESET_B(net75),
    .D(_0057_),
    .Q(\ayayayayayaya.b[25] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_1 _3487_ (.RESET_B(net74),
    .D(_0058_),
    .Q(\ayayayayayaya.b[26] ),
    .CLK(clknet_4_9_0_clk));
 sg13g2_dfrbpq_2 _3488_ (.RESET_B(net73),
    .D(_0059_),
    .Q(\ayayayayayaya.b[27] ),
    .CLK(clknet_4_14_0_clk));
 sg13g2_dfrbpq_2 _3489_ (.RESET_B(net72),
    .D(_0060_),
    .Q(\ayayayayayaya.b[28] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _3490_ (.RESET_B(net71),
    .D(_0061_),
    .Q(\ayayayayayaya.b[29] ),
    .CLK(clknet_4_12_0_clk));
 sg13g2_dfrbpq_2 _3491_ (.RESET_B(net70),
    .D(_0062_),
    .Q(\ayayayayayaya.b[30] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_dfrbpq_2 _3492_ (.RESET_B(net69),
    .D(_0063_),
    .Q(\ayayayayayaya.b[31] ),
    .CLK(clknet_4_13_0_clk));
 sg13g2_tiehi _3482__15 (.L_HI(net15));
 sg13g2_tiehi _3481__16 (.L_HI(net16));
 sg13g2_tiehi _3480__17 (.L_HI(net17));
 sg13g2_tiehi _3479__18 (.L_HI(net18));
 sg13g2_tiehi _3478__19 (.L_HI(net19));
 sg13g2_tiehi _3477__20 (.L_HI(net20));
 sg13g2_tiehi _3476__21 (.L_HI(net21));
 sg13g2_tiehi _3475__22 (.L_HI(net22));
 sg13g2_tiehi _3474__23 (.L_HI(net23));
 sg13g2_tiehi _3473__24 (.L_HI(net24));
 sg13g2_tiehi _3472__25 (.L_HI(net25));
 sg13g2_tiehi _3471__26 (.L_HI(net26));
 sg13g2_tiehi _3470__27 (.L_HI(net27));
 sg13g2_tiehi _3469__28 (.L_HI(net28));
 sg13g2_tiehi _3468__29 (.L_HI(net29));
 sg13g2_tiehi _3467__30 (.L_HI(net30));
 sg13g2_tiehi _3466__31 (.L_HI(net31));
 sg13g2_tiehi _3465__32 (.L_HI(net32));
 sg13g2_tiehi _3464__33 (.L_HI(net33));
 sg13g2_tiehi _3463__34 (.L_HI(net34));
 sg13g2_tiehi _3462__35 (.L_HI(net35));
 sg13g2_tiehi _3461__36 (.L_HI(net36));
 sg13g2_tiehi _3460__37 (.L_HI(net37));
 sg13g2_tiehi _3459__38 (.L_HI(net38));
 sg13g2_tiehi _3458__39 (.L_HI(net39));
 sg13g2_tiehi _3457__40 (.L_HI(net40));
 sg13g2_tiehi _3456__41 (.L_HI(net41));
 sg13g2_tiehi _3455__42 (.L_HI(net42));
 sg13g2_tiehi _3454__43 (.L_HI(net43));
 sg13g2_tiehi _3453__44 (.L_HI(net44));
 sg13g2_tiehi _3452__45 (.L_HI(net45));
 sg13g2_tiehi _3451__46 (.L_HI(net46));
 sg13g2_tiehi _3450__47 (.L_HI(net47));
 sg13g2_tiehi _3449__48 (.L_HI(net48));
 sg13g2_tiehi _3448__49 (.L_HI(net49));
 sg13g2_tiehi _3447__50 (.L_HI(net50));
 sg13g2_tiehi _3446__51 (.L_HI(net51));
 sg13g2_tiehi _3445__52 (.L_HI(net52));
 sg13g2_tiehi _3444__53 (.L_HI(net53));
 sg13g2_tiehi _3443__54 (.L_HI(net54));
 sg13g2_tiehi _3442__55 (.L_HI(net55));
 sg13g2_tiehi _3441__56 (.L_HI(net56));
 sg13g2_tiehi _3440__57 (.L_HI(net57));
 sg13g2_tiehi _3439__58 (.L_HI(net58));
 sg13g2_tiehi _3438__59 (.L_HI(net59));
 sg13g2_tiehi _3437__60 (.L_HI(net60));
 sg13g2_tiehi _3436__61 (.L_HI(net61));
 sg13g2_tiehi _3435__62 (.L_HI(net62));
 sg13g2_tiehi _3434__63 (.L_HI(net63));
 sg13g2_tiehi _3433__64 (.L_HI(net64));
 sg13g2_tiehi _3432__65 (.L_HI(net65));
 sg13g2_tiehi _3431__66 (.L_HI(net66));
 sg13g2_tiehi _3430__67 (.L_HI(net67));
 sg13g2_tiehi _3429__68 (.L_HI(net68));
 sg13g2_tiehi _3492__69 (.L_HI(net69));
 sg13g2_tiehi _3491__70 (.L_HI(net70));
 sg13g2_tiehi _3490__71 (.L_HI(net71));
 sg13g2_tiehi _3489__72 (.L_HI(net72));
 sg13g2_tiehi _3488__73 (.L_HI(net73));
 sg13g2_tiehi _3487__74 (.L_HI(net74));
 sg13g2_tiehi _3486__75 (.L_HI(net75));
 sg13g2_tiehi _3485__76 (.L_HI(net76));
 sg13g2_tiehi _3484__77 (.L_HI(net77));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_buf_1 _3557_ (.A(uio_oe[7]),
    .X(uio_oe[0]));
 sg13g2_buf_1 _3558_ (.A(uio_oe[7]),
    .X(uio_oe[1]));
 sg13g2_buf_1 _3559_ (.A(uio_oe[7]),
    .X(uio_oe[2]));
 sg13g2_buf_1 _3560_ (.A(uio_oe[7]),
    .X(uio_oe[3]));
 sg13g2_buf_1 _3561_ (.A(uio_oe[7]),
    .X(uio_oe[4]));
 sg13g2_buf_1 _3562_ (.A(uio_oe[7]),
    .X(uio_oe[5]));
 sg13g2_buf_1 _3563_ (.A(uio_oe[7]),
    .X(uio_oe[6]));
 sg13g2_buf_1 _3564_ (.A(uio_out[0]),
    .X(uo_out[0]));
 sg13g2_buf_1 _3565_ (.A(uio_out[1]),
    .X(uo_out[1]));
 sg13g2_buf_1 _3566_ (.A(uio_out[2]),
    .X(uo_out[2]));
 sg13g2_buf_1 _3567_ (.A(uio_out[3]),
    .X(uo_out[3]));
 sg13g2_buf_1 _3568_ (.A(uio_out[4]),
    .X(uo_out[4]));
 sg13g2_buf_1 _3569_ (.A(uio_out[5]),
    .X(uo_out[5]));
 sg13g2_buf_1 _3570_ (.A(uio_out[6]),
    .X(uo_out[6]));
 sg13g2_buf_1 _3571_ (.A(uio_out[7]),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout578 (.A(_0855_),
    .X(net578));
 sg13g2_buf_2 fanout579 (.A(_0855_),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(_0844_),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(_0844_),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(_0834_),
    .X(net582));
 sg13g2_buf_8 fanout583 (.A(_0834_),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584));
 sg13g2_buf_8 fanout585 (.A(_0824_),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(_0821_),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(_0815_),
    .X(net587));
 sg13g2_buf_8 fanout588 (.A(_0812_),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net590),
    .X(net589));
 sg13g2_buf_8 fanout590 (.A(_0188_),
    .X(net590));
 sg13g2_buf_8 fanout591 (.A(net592),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(_0112_),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net597),
    .X(net593));
 sg13g2_buf_1 fanout594 (.A(net597),
    .X(net594));
 sg13g2_buf_2 fanout595 (.A(net596),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_2 fanout597 (.A(_1370_),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(_0872_),
    .X(net598));
 sg13g2_buf_1 fanout599 (.A(_0872_),
    .X(net599));
 sg13g2_buf_2 fanout600 (.A(net601),
    .X(net600));
 sg13g2_buf_8 fanout601 (.A(_0872_),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net603),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(_1424_),
    .X(net603));
 sg13g2_buf_8 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(_1412_),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(_1411_),
    .X(net606));
 sg13g2_buf_1 fanout607 (.A(_1411_),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(_1410_),
    .X(net609));
 sg13g2_buf_8 fanout610 (.A(_1410_),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(net612),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_1 fanout613 (.A(_1408_),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_8 fanout615 (.A(_1408_),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net617),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net618),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(_1404_),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(_1404_),
    .X(net619));
 sg13g2_buf_1 fanout620 (.A(_1404_),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net622),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(_1402_),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(net625),
    .X(net623));
 sg13g2_buf_1 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(_1402_),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(net628),
    .X(net626));
 sg13g2_buf_1 fanout627 (.A(net628),
    .X(net627));
 sg13g2_buf_2 fanout628 (.A(net629),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(_0868_),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(_0868_),
    .X(net630));
 sg13g2_buf_1 fanout631 (.A(net632),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(_0868_),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net635),
    .X(net633));
 sg13g2_buf_2 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net639),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net639),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(net639),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(_0867_),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(net642),
    .X(net640));
 sg13g2_buf_1 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(_0866_),
    .X(net642));
 sg13g2_buf_2 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(_0866_),
    .X(net644));
 sg13g2_buf_8 fanout645 (.A(_0866_),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(net648),
    .X(net646));
 sg13g2_buf_1 fanout647 (.A(net648),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(net653),
    .X(net648));
 sg13g2_buf_2 fanout649 (.A(net650),
    .X(net649));
 sg13g2_buf_1 fanout650 (.A(net653),
    .X(net650));
 sg13g2_buf_2 fanout651 (.A(net652),
    .X(net651));
 sg13g2_buf_1 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_1 fanout653 (.A(_0865_),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_2 fanout655 (.A(_0864_),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(net657),
    .X(net656));
 sg13g2_buf_2 fanout657 (.A(net658),
    .X(net657));
 sg13g2_buf_8 fanout658 (.A(_0864_),
    .X(net658));
 sg13g2_buf_8 fanout659 (.A(net660),
    .X(net659));
 sg13g2_buf_8 fanout660 (.A(_0863_),
    .X(net660));
 sg13g2_buf_8 fanout661 (.A(net662),
    .X(net661));
 sg13g2_buf_1 fanout662 (.A(net663),
    .X(net662));
 sg13g2_buf_8 fanout663 (.A(_0863_),
    .X(net663));
 sg13g2_buf_8 fanout664 (.A(net665),
    .X(net664));
 sg13g2_buf_2 fanout665 (.A(_0858_),
    .X(net665));
 sg13g2_buf_2 fanout666 (.A(net667),
    .X(net666));
 sg13g2_buf_1 fanout667 (.A(net668),
    .X(net667));
 sg13g2_buf_8 fanout668 (.A(_0858_),
    .X(net668));
 sg13g2_buf_8 fanout669 (.A(net673),
    .X(net669));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670));
 sg13g2_buf_2 fanout671 (.A(net672),
    .X(net671));
 sg13g2_buf_2 fanout672 (.A(net673),
    .X(net672));
 sg13g2_buf_1 fanout673 (.A(_0851_),
    .X(net673));
 sg13g2_buf_8 fanout674 (.A(net675),
    .X(net674));
 sg13g2_buf_1 fanout675 (.A(net678),
    .X(net675));
 sg13g2_buf_8 fanout676 (.A(net677),
    .X(net676));
 sg13g2_buf_8 fanout677 (.A(net678),
    .X(net677));
 sg13g2_buf_1 fanout678 (.A(_0845_),
    .X(net678));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679));
 sg13g2_buf_8 fanout680 (.A(net681),
    .X(net680));
 sg13g2_buf_8 fanout681 (.A(_0839_),
    .X(net681));
 sg13g2_buf_2 fanout682 (.A(net684),
    .X(net682));
 sg13g2_buf_1 fanout683 (.A(net684),
    .X(net683));
 sg13g2_buf_1 fanout684 (.A(net685),
    .X(net684));
 sg13g2_buf_8 fanout685 (.A(_0832_),
    .X(net685));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686));
 sg13g2_buf_2 fanout687 (.A(net688),
    .X(net687));
 sg13g2_buf_8 fanout688 (.A(_0826_),
    .X(net688));
 sg13g2_buf_2 fanout689 (.A(net690),
    .X(net689));
 sg13g2_buf_1 fanout690 (.A(net691),
    .X(net690));
 sg13g2_buf_1 fanout691 (.A(_0823_),
    .X(net691));
 sg13g2_buf_8 fanout692 (.A(_0823_),
    .X(net692));
 sg13g2_buf_8 fanout693 (.A(net695),
    .X(net693));
 sg13g2_buf_1 fanout694 (.A(net695),
    .X(net694));
 sg13g2_buf_1 fanout695 (.A(net696),
    .X(net695));
 sg13g2_buf_1 fanout696 (.A(_0818_),
    .X(net696));
 sg13g2_buf_8 fanout697 (.A(net698),
    .X(net697));
 sg13g2_buf_8 fanout698 (.A(_0813_),
    .X(net698));
 sg13g2_buf_8 fanout699 (.A(net700),
    .X(net699));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700));
 sg13g2_buf_1 fanout701 (.A(_0810_),
    .X(net701));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702));
 sg13g2_buf_8 fanout703 (.A(_0806_),
    .X(net703));
 sg13g2_buf_8 fanout704 (.A(net705),
    .X(net704));
 sg13g2_buf_8 fanout705 (.A(_0795_),
    .X(net705));
 sg13g2_buf_8 fanout706 (.A(net707),
    .X(net706));
 sg13g2_buf_8 fanout707 (.A(_0784_),
    .X(net707));
 sg13g2_buf_8 fanout708 (.A(_0773_),
    .X(net708));
 sg13g2_buf_1 fanout709 (.A(_0773_),
    .X(net709));
 sg13g2_buf_8 fanout710 (.A(_0762_),
    .X(net710));
 sg13g2_buf_8 fanout711 (.A(_0751_),
    .X(net711));
 sg13g2_buf_1 fanout712 (.A(_0751_),
    .X(net712));
 sg13g2_buf_8 fanout713 (.A(_0740_),
    .X(net713));
 sg13g2_buf_8 fanout714 (.A(_0730_),
    .X(net714));
 sg13g2_buf_8 fanout715 (.A(_0719_),
    .X(net715));
 sg13g2_buf_8 fanout716 (.A(net116),
    .X(net716));
 sg13g2_buf_8 fanout717 (.A(net118),
    .X(net717));
 sg13g2_buf_8 fanout718 (.A(\ayayayayayaya.b[24] ),
    .X(net718));
 sg13g2_buf_8 fanout719 (.A(net720),
    .X(net719));
 sg13g2_buf_8 fanout720 (.A(\ayayayayayaya.b[23] ),
    .X(net720));
 sg13g2_buf_8 fanout721 (.A(\ayayayayayaya.b[22] ),
    .X(net721));
 sg13g2_buf_8 fanout722 (.A(net724),
    .X(net722));
 sg13g2_buf_1 fanout723 (.A(net724),
    .X(net723));
 sg13g2_buf_8 fanout724 (.A(\ayayayayayaya.b[21] ),
    .X(net724));
 sg13g2_buf_2 fanout725 (.A(net726),
    .X(net725));
 sg13g2_buf_8 fanout726 (.A(net117),
    .X(net726));
 sg13g2_buf_8 fanout727 (.A(net728),
    .X(net727));
 sg13g2_buf_8 fanout728 (.A(\ayayayayayaya.b[19] ),
    .X(net728));
 sg13g2_buf_2 fanout729 (.A(net730),
    .X(net729));
 sg13g2_buf_8 fanout730 (.A(\ayayayayayaya.b[18] ),
    .X(net730));
 sg13g2_buf_2 fanout731 (.A(net732),
    .X(net731));
 sg13g2_buf_1 fanout732 (.A(net733),
    .X(net732));
 sg13g2_buf_1 fanout733 (.A(net734),
    .X(net733));
 sg13g2_buf_2 fanout734 (.A(\ayayayayayaya.b[17] ),
    .X(net734));
 sg13g2_buf_2 fanout735 (.A(net736),
    .X(net735));
 sg13g2_buf_1 fanout736 (.A(net737),
    .X(net736));
 sg13g2_buf_8 fanout737 (.A(\ayayayayayaya.b[16] ),
    .X(net737));
 sg13g2_buf_2 fanout738 (.A(net739),
    .X(net738));
 sg13g2_buf_1 fanout739 (.A(net740),
    .X(net739));
 sg13g2_buf_1 fanout740 (.A(net741),
    .X(net740));
 sg13g2_buf_8 fanout741 (.A(\ayayayayayaya.b[15] ),
    .X(net741));
 sg13g2_buf_2 fanout742 (.A(net743),
    .X(net742));
 sg13g2_buf_1 fanout743 (.A(net744),
    .X(net743));
 sg13g2_buf_1 fanout744 (.A(\ayayayayayaya.b[14] ),
    .X(net744));
 sg13g2_buf_8 fanout745 (.A(\ayayayayayaya.b[14] ),
    .X(net745));
 sg13g2_buf_2 fanout746 (.A(net747),
    .X(net746));
 sg13g2_buf_1 fanout747 (.A(net748),
    .X(net747));
 sg13g2_buf_8 fanout748 (.A(\ayayayayayaya.b[13] ),
    .X(net748));
 sg13g2_buf_8 fanout749 (.A(\ayayayayayaya.b[12] ),
    .X(net749));
 sg13g2_buf_2 fanout750 (.A(net752),
    .X(net750));
 sg13g2_buf_1 fanout751 (.A(net752),
    .X(net751));
 sg13g2_buf_1 fanout752 (.A(\ayayayayayaya.b[12] ),
    .X(net752));
 sg13g2_buf_8 fanout753 (.A(net754),
    .X(net753));
 sg13g2_buf_8 fanout754 (.A(\ayayayayayaya.b[11] ),
    .X(net754));
 sg13g2_buf_2 fanout755 (.A(net756),
    .X(net755));
 sg13g2_buf_8 fanout756 (.A(\ayayayayayaya.b[11] ),
    .X(net756));
 sg13g2_buf_2 fanout757 (.A(net758),
    .X(net757));
 sg13g2_buf_1 fanout758 (.A(net759),
    .X(net758));
 sg13g2_buf_1 fanout759 (.A(net762),
    .X(net759));
 sg13g2_buf_8 fanout760 (.A(net761),
    .X(net760));
 sg13g2_buf_8 fanout761 (.A(net762),
    .X(net761));
 sg13g2_buf_8 fanout762 (.A(\ayayayayayaya.b[10] ),
    .X(net762));
 sg13g2_buf_8 fanout763 (.A(net767),
    .X(net763));
 sg13g2_buf_1 fanout764 (.A(net767),
    .X(net764));
 sg13g2_buf_8 fanout765 (.A(net766),
    .X(net765));
 sg13g2_buf_8 fanout766 (.A(net767),
    .X(net766));
 sg13g2_buf_8 fanout767 (.A(\ayayayayayaya.b[9] ),
    .X(net767));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768));
 sg13g2_buf_8 fanout769 (.A(net773),
    .X(net769));
 sg13g2_buf_8 fanout770 (.A(net772),
    .X(net770));
 sg13g2_buf_1 fanout771 (.A(net772),
    .X(net771));
 sg13g2_buf_8 fanout772 (.A(net773),
    .X(net772));
 sg13g2_buf_8 fanout773 (.A(\ayayayayayaya.b[8] ),
    .X(net773));
 sg13g2_buf_8 fanout774 (.A(net775),
    .X(net774));
 sg13g2_buf_2 fanout775 (.A(net779),
    .X(net775));
 sg13g2_buf_2 fanout776 (.A(net777),
    .X(net776));
 sg13g2_buf_1 fanout777 (.A(net778),
    .X(net777));
 sg13g2_buf_1 fanout778 (.A(net779),
    .X(net778));
 sg13g2_buf_8 fanout779 (.A(\ayayayayayaya.b[7] ),
    .X(net779));
 sg13g2_buf_8 fanout780 (.A(net781),
    .X(net780));
 sg13g2_buf_8 fanout781 (.A(net785),
    .X(net781));
 sg13g2_buf_8 fanout782 (.A(net783),
    .X(net782));
 sg13g2_buf_8 fanout783 (.A(net784),
    .X(net783));
 sg13g2_buf_8 fanout784 (.A(net785),
    .X(net784));
 sg13g2_buf_8 fanout785 (.A(\ayayayayayaya.b[6] ),
    .X(net785));
 sg13g2_buf_8 fanout786 (.A(net787),
    .X(net786));
 sg13g2_buf_8 fanout787 (.A(net788),
    .X(net787));
 sg13g2_buf_8 fanout788 (.A(net792),
    .X(net788));
 sg13g2_buf_8 fanout789 (.A(net792),
    .X(net789));
 sg13g2_buf_8 fanout790 (.A(net791),
    .X(net790));
 sg13g2_buf_2 fanout791 (.A(net792),
    .X(net791));
 sg13g2_buf_8 fanout792 (.A(\ayayayayayaya.b[5] ),
    .X(net792));
 sg13g2_buf_8 fanout793 (.A(net794),
    .X(net793));
 sg13g2_buf_8 fanout794 (.A(net795),
    .X(net794));
 sg13g2_buf_2 fanout795 (.A(net799),
    .X(net795));
 sg13g2_buf_2 fanout796 (.A(net799),
    .X(net796));
 sg13g2_buf_1 fanout797 (.A(net799),
    .X(net797));
 sg13g2_buf_2 fanout798 (.A(net799),
    .X(net798));
 sg13g2_buf_1 fanout799 (.A(\ayayayayayaya.b[4] ),
    .X(net799));
 sg13g2_buf_8 fanout800 (.A(net802),
    .X(net800));
 sg13g2_buf_1 fanout801 (.A(net802),
    .X(net801));
 sg13g2_buf_8 fanout802 (.A(\ayayayayayaya.b[3] ),
    .X(net802));
 sg13g2_buf_8 fanout803 (.A(net806),
    .X(net803));
 sg13g2_buf_2 fanout804 (.A(net806),
    .X(net804));
 sg13g2_buf_1 fanout805 (.A(net806),
    .X(net805));
 sg13g2_buf_2 fanout806 (.A(\ayayayayayaya.b[3] ),
    .X(net806));
 sg13g2_buf_8 fanout807 (.A(net809),
    .X(net807));
 sg13g2_buf_8 fanout808 (.A(net809),
    .X(net808));
 sg13g2_buf_8 fanout809 (.A(\ayayayayayaya.b[2] ),
    .X(net809));
 sg13g2_buf_2 fanout810 (.A(net812),
    .X(net810));
 sg13g2_buf_1 fanout811 (.A(net812),
    .X(net811));
 sg13g2_buf_2 fanout812 (.A(net813),
    .X(net812));
 sg13g2_buf_1 fanout813 (.A(\ayayayayayaya.b[2] ),
    .X(net813));
 sg13g2_buf_8 fanout814 (.A(net817),
    .X(net814));
 sg13g2_buf_1 fanout815 (.A(net817),
    .X(net815));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816));
 sg13g2_buf_8 fanout817 (.A(net821),
    .X(net817));
 sg13g2_buf_2 fanout818 (.A(net820),
    .X(net818));
 sg13g2_buf_1 fanout819 (.A(net820),
    .X(net819));
 sg13g2_buf_1 fanout820 (.A(net821),
    .X(net820));
 sg13g2_buf_1 fanout821 (.A(\ayayayayayaya.b[1] ),
    .X(net821));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822));
 sg13g2_buf_2 fanout823 (.A(net113),
    .X(net823));
 sg13g2_buf_8 fanout824 (.A(\a[15] ),
    .X(net824));
 sg13g2_buf_8 fanout825 (.A(\a[8] ),
    .X(net825));
 sg13g2_buf_8 fanout826 (.A(\a[7] ),
    .X(net826));
 sg13g2_buf_8 fanout827 (.A(net828),
    .X(net827));
 sg13g2_buf_2 fanout828 (.A(\a[0] ),
    .X(net828));
 sg13g2_buf_8 fanout829 (.A(net115),
    .X(net829));
 sg13g2_buf_8 fanout830 (.A(net114),
    .X(net830));
 sg13g2_buf_1 fanout831 (.A(\a[16] ),
    .X(net831));
 sg13g2_buf_8 fanout832 (.A(net833),
    .X(net832));
 sg13g2_buf_8 fanout833 (.A(_1417_),
    .X(net833));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834));
 sg13g2_buf_8 fanout835 (.A(net836),
    .X(net835));
 sg13g2_buf_2 fanout836 (.A(_1417_),
    .X(net836));
 sg13g2_buf_8 fanout837 (.A(_1416_),
    .X(net837));
 sg13g2_buf_8 fanout838 (.A(_1406_),
    .X(net838));
 sg13g2_buf_8 fanout839 (.A(net842),
    .X(net839));
 sg13g2_buf_2 fanout840 (.A(net842),
    .X(net840));
 sg13g2_buf_8 fanout841 (.A(net842),
    .X(net841));
 sg13g2_buf_8 fanout842 (.A(ui_in[3]),
    .X(net842));
 sg13g2_buf_8 fanout843 (.A(net844),
    .X(net843));
 sg13g2_buf_8 fanout844 (.A(ui_in[1]),
    .X(net844));
 sg13g2_buf_8 fanout845 (.A(net846),
    .X(net845));
 sg13g2_buf_8 fanout846 (.A(ui_in[0]),
    .X(net846));
 sg13g2_buf_2 fanout847 (.A(ui_in[0]),
    .X(net847));
 sg13g2_buf_8 fanout848 (.A(net849),
    .X(net848));
 sg13g2_buf_8 fanout849 (.A(ui_in[0]),
    .X(net849));
 sg13g2_buf_2 input1 (.A(ui_in[2]),
    .X(net1));
 sg13g2_buf_2 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_2 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_2 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_2 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_2 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_2 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_2 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_2 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_2 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_2 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_buf_2 input13 (.A(uio_in[7]),
    .X(net13));
 sg13g2_tiehi _3483__14 (.L_HI(net14));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_4_0_0_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_4_1_0_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_4_2_0_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_4_3_0_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_4_4_0_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_4_5_0_clk));
 sg13g2_buf_1 clkload6 (.A(clknet_4_7_0_clk));
 sg13g2_buf_1 clkload7 (.A(clknet_4_8_0_clk));
 sg13g2_buf_1 clkload8 (.A(clknet_4_9_0_clk));
 sg13g2_buf_1 clkload9 (.A(clknet_4_10_0_clk));
 sg13g2_buf_1 clkload10 (.A(clknet_4_11_0_clk));
 sg13g2_buf_1 clkload11 (.A(clknet_4_15_0_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\a[0] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold2 (.A(\a[7] ),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold3 (.A(\a[8] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold4 (.A(\a[1] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold5 (.A(\a[5] ),
    .X(net82));
 sg13g2_dlygate4sd3_1 hold6 (.A(\a[15] ),
    .X(net83));
 sg13g2_dlygate4sd3_1 hold7 (.A(\a[26] ),
    .X(net84));
 sg13g2_dlygate4sd3_1 hold8 (.A(\ayayayayayaya.b[30] ),
    .X(net85));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ayayayayayaya.b[31] ),
    .X(net86));
 sg13g2_dlygate4sd3_1 hold10 (.A(\ayayayayayaya.b[28] ),
    .X(net87));
 sg13g2_dlygate4sd3_1 hold11 (.A(\a[30] ),
    .X(net88));
 sg13g2_dlygate4sd3_1 hold12 (.A(\a[27] ),
    .X(net89));
 sg13g2_dlygate4sd3_1 hold13 (.A(\a[25] ),
    .X(net90));
 sg13g2_dlygate4sd3_1 hold14 (.A(\ayayayayayaya.b[29] ),
    .X(net91));
 sg13g2_dlygate4sd3_1 hold15 (.A(\a[24] ),
    .X(net92));
 sg13g2_dlygate4sd3_1 hold16 (.A(\a[10] ),
    .X(net93));
 sg13g2_dlygate4sd3_1 hold17 (.A(\a[11] ),
    .X(net94));
 sg13g2_dlygate4sd3_1 hold18 (.A(\a[2] ),
    .X(net95));
 sg13g2_dlygate4sd3_1 hold19 (.A(\a[29] ),
    .X(net96));
 sg13g2_dlygate4sd3_1 hold20 (.A(\a[19] ),
    .X(net97));
 sg13g2_dlygate4sd3_1 hold21 (.A(\a[21] ),
    .X(net98));
 sg13g2_dlygate4sd3_1 hold22 (.A(\a[14] ),
    .X(net99));
 sg13g2_dlygate4sd3_1 hold23 (.A(\a[3] ),
    .X(net100));
 sg13g2_dlygate4sd3_1 hold24 (.A(\a[9] ),
    .X(net101));
 sg13g2_dlygate4sd3_1 hold25 (.A(\a[28] ),
    .X(net102));
 sg13g2_dlygate4sd3_1 hold26 (.A(\a[6] ),
    .X(net103));
 sg13g2_dlygate4sd3_1 hold27 (.A(\a[13] ),
    .X(net104));
 sg13g2_dlygate4sd3_1 hold28 (.A(\a[4] ),
    .X(net105));
 sg13g2_dlygate4sd3_1 hold29 (.A(\a[23] ),
    .X(net106));
 sg13g2_dlygate4sd3_1 hold30 (.A(\a[17] ),
    .X(net107));
 sg13g2_dlygate4sd3_1 hold31 (.A(\a[12] ),
    .X(net108));
 sg13g2_dlygate4sd3_1 hold32 (.A(\a[22] ),
    .X(net109));
 sg13g2_dlygate4sd3_1 hold33 (.A(\a[20] ),
    .X(net110));
 sg13g2_dlygate4sd3_1 hold34 (.A(\ayayayayayaya.b[27] ),
    .X(net111));
 sg13g2_dlygate4sd3_1 hold35 (.A(\a[18] ),
    .X(net112));
 sg13g2_dlygate4sd3_1 hold36 (.A(\ayayayayayaya.b[0] ),
    .X(net113));
 sg13g2_dlygate4sd3_1 hold37 (.A(\a[16] ),
    .X(net114));
 sg13g2_dlygate4sd3_1 hold38 (.A(\a[31] ),
    .X(net115));
 sg13g2_dlygate4sd3_1 hold39 (.A(\ayayayayayaya.b[26] ),
    .X(net116));
 sg13g2_dlygate4sd3_1 hold40 (.A(\ayayayayayaya.b[20] ),
    .X(net117));
 sg13g2_dlygate4sd3_1 hold41 (.A(\ayayayayayaya.b[25] ),
    .X(net118));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_39 ();
 sg13g2_fill_2 FILLER_0_46 ();
 sg13g2_fill_1 FILLER_0_48 ();
 sg13g2_fill_2 FILLER_0_73 ();
 sg13g2_fill_1 FILLER_0_100 ();
 sg13g2_fill_2 FILLER_0_125 ();
 sg13g2_fill_2 FILLER_0_155 ();
 sg13g2_fill_1 FILLER_0_157 ();
 sg13g2_fill_2 FILLER_0_167 ();
 sg13g2_fill_1 FILLER_0_169 ();
 sg13g2_fill_1 FILLER_0_187 ();
 sg13g2_decap_8 FILLER_0_206 ();
 sg13g2_fill_2 FILLER_0_213 ();
 sg13g2_fill_1 FILLER_0_232 ();
 sg13g2_decap_4 FILLER_0_247 ();
 sg13g2_decap_8 FILLER_0_256 ();
 sg13g2_fill_2 FILLER_0_263 ();
 sg13g2_fill_1 FILLER_0_265 ();
 sg13g2_decap_8 FILLER_0_271 ();
 sg13g2_decap_4 FILLER_0_282 ();
 sg13g2_fill_1 FILLER_0_286 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_fill_2 FILLER_0_297 ();
 sg13g2_decap_4 FILLER_0_304 ();
 sg13g2_fill_1 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_324 ();
 sg13g2_fill_1 FILLER_0_331 ();
 sg13g2_decap_8 FILLER_0_375 ();
 sg13g2_decap_8 FILLER_0_382 ();
 sg13g2_decap_8 FILLER_0_389 ();
 sg13g2_decap_8 FILLER_0_396 ();
 sg13g2_decap_4 FILLER_0_403 ();
 sg13g2_fill_2 FILLER_0_407 ();
 sg13g2_fill_2 FILLER_1_0 ();
 sg13g2_fill_1 FILLER_1_2 ();
 sg13g2_decap_8 FILLER_1_11 ();
 sg13g2_decap_8 FILLER_1_18 ();
 sg13g2_fill_1 FILLER_1_25 ();
 sg13g2_fill_2 FILLER_1_46 ();
 sg13g2_fill_1 FILLER_1_48 ();
 sg13g2_fill_2 FILLER_1_78 ();
 sg13g2_fill_1 FILLER_1_80 ();
 sg13g2_fill_1 FILLER_1_94 ();
 sg13g2_fill_2 FILLER_1_105 ();
 sg13g2_fill_1 FILLER_1_107 ();
 sg13g2_fill_2 FILLER_1_123 ();
 sg13g2_fill_2 FILLER_1_130 ();
 sg13g2_fill_2 FILLER_1_156 ();
 sg13g2_fill_1 FILLER_1_158 ();
 sg13g2_fill_2 FILLER_1_207 ();
 sg13g2_fill_1 FILLER_1_209 ();
 sg13g2_fill_2 FILLER_1_254 ();
 sg13g2_fill_2 FILLER_1_265 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_fill_2 FILLER_1_329 ();
 sg13g2_fill_1 FILLER_1_374 ();
 sg13g2_decap_8 FILLER_1_388 ();
 sg13g2_decap_8 FILLER_1_395 ();
 sg13g2_decap_8 FILLER_1_402 ();
 sg13g2_fill_2 FILLER_2_0 ();
 sg13g2_fill_1 FILLER_2_2 ();
 sg13g2_fill_1 FILLER_2_11 ();
 sg13g2_fill_2 FILLER_2_16 ();
 sg13g2_fill_1 FILLER_2_18 ();
 sg13g2_fill_2 FILLER_2_39 ();
 sg13g2_fill_1 FILLER_2_41 ();
 sg13g2_fill_2 FILLER_2_77 ();
 sg13g2_fill_1 FILLER_2_79 ();
 sg13g2_fill_1 FILLER_2_105 ();
 sg13g2_fill_1 FILLER_2_120 ();
 sg13g2_fill_1 FILLER_2_131 ();
 sg13g2_fill_2 FILLER_2_142 ();
 sg13g2_fill_1 FILLER_2_164 ();
 sg13g2_fill_2 FILLER_2_170 ();
 sg13g2_fill_1 FILLER_2_172 ();
 sg13g2_fill_2 FILLER_2_183 ();
 sg13g2_decap_4 FILLER_2_209 ();
 sg13g2_fill_1 FILLER_2_213 ();
 sg13g2_decap_4 FILLER_2_229 ();
 sg13g2_fill_1 FILLER_2_233 ();
 sg13g2_decap_4 FILLER_2_278 ();
 sg13g2_fill_2 FILLER_2_302 ();
 sg13g2_fill_2 FILLER_2_319 ();
 sg13g2_fill_1 FILLER_2_321 ();
 sg13g2_fill_2 FILLER_2_332 ();
 sg13g2_fill_2 FILLER_2_369 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_4 FILLER_2_403 ();
 sg13g2_fill_2 FILLER_2_407 ();
 sg13g2_fill_1 FILLER_3_0 ();
 sg13g2_decap_4 FILLER_3_45 ();
 sg13g2_fill_1 FILLER_3_49 ();
 sg13g2_decap_4 FILLER_3_74 ();
 sg13g2_fill_2 FILLER_3_78 ();
 sg13g2_fill_1 FILLER_3_100 ();
 sg13g2_fill_2 FILLER_3_181 ();
 sg13g2_fill_1 FILLER_3_188 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_2 FILLER_3_223 ();
 sg13g2_fill_2 FILLER_3_235 ();
 sg13g2_fill_1 FILLER_3_251 ();
 sg13g2_fill_1 FILLER_3_257 ();
 sg13g2_fill_2 FILLER_3_263 ();
 sg13g2_fill_1 FILLER_3_265 ();
 sg13g2_decap_4 FILLER_3_300 ();
 sg13g2_fill_2 FILLER_3_324 ();
 sg13g2_fill_1 FILLER_3_326 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_fill_2 FILLER_3_406 ();
 sg13g2_fill_1 FILLER_3_408 ();
 sg13g2_fill_2 FILLER_4_0 ();
 sg13g2_fill_1 FILLER_4_2 ();
 sg13g2_fill_2 FILLER_4_16 ();
 sg13g2_decap_4 FILLER_4_58 ();
 sg13g2_fill_1 FILLER_4_79 ();
 sg13g2_fill_1 FILLER_4_95 ();
 sg13g2_fill_2 FILLER_4_121 ();
 sg13g2_fill_2 FILLER_4_164 ();
 sg13g2_fill_1 FILLER_4_178 ();
 sg13g2_fill_2 FILLER_4_204 ();
 sg13g2_fill_1 FILLER_4_206 ();
 sg13g2_fill_2 FILLER_4_217 ();
 sg13g2_fill_1 FILLER_4_219 ();
 sg13g2_fill_1 FILLER_4_238 ();
 sg13g2_fill_1 FILLER_4_267 ();
 sg13g2_fill_2 FILLER_4_313 ();
 sg13g2_fill_1 FILLER_4_315 ();
 sg13g2_fill_2 FILLER_4_356 ();
 sg13g2_fill_1 FILLER_4_358 ();
 sg13g2_fill_2 FILLER_5_4 ();
 sg13g2_fill_1 FILLER_5_6 ();
 sg13g2_fill_2 FILLER_5_30 ();
 sg13g2_fill_1 FILLER_5_52 ();
 sg13g2_fill_2 FILLER_5_63 ();
 sg13g2_fill_1 FILLER_5_65 ();
 sg13g2_fill_2 FILLER_5_75 ();
 sg13g2_fill_1 FILLER_5_115 ();
 sg13g2_fill_1 FILLER_5_134 ();
 sg13g2_fill_2 FILLER_5_166 ();
 sg13g2_decap_4 FILLER_5_201 ();
 sg13g2_fill_1 FILLER_5_205 ();
 sg13g2_decap_8 FILLER_5_216 ();
 sg13g2_fill_1 FILLER_5_223 ();
 sg13g2_fill_2 FILLER_5_255 ();
 sg13g2_fill_2 FILLER_5_262 ();
 sg13g2_fill_1 FILLER_5_264 ();
 sg13g2_fill_1 FILLER_5_270 ();
 sg13g2_decap_4 FILLER_5_296 ();
 sg13g2_fill_1 FILLER_5_320 ();
 sg13g2_decap_4 FILLER_5_336 ();
 sg13g2_fill_2 FILLER_5_353 ();
 sg13g2_fill_2 FILLER_5_365 ();
 sg13g2_decap_8 FILLER_6_40 ();
 sg13g2_fill_1 FILLER_6_47 ();
 sg13g2_decap_4 FILLER_6_58 ();
 sg13g2_fill_2 FILLER_6_62 ();
 sg13g2_fill_1 FILLER_6_79 ();
 sg13g2_fill_2 FILLER_6_90 ();
 sg13g2_fill_1 FILLER_6_92 ();
 sg13g2_fill_2 FILLER_6_123 ();
 sg13g2_fill_1 FILLER_6_133 ();
 sg13g2_fill_2 FILLER_6_152 ();
 sg13g2_fill_1 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_174 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_fill_1 FILLER_6_200 ();
 sg13g2_fill_1 FILLER_6_211 ();
 sg13g2_fill_2 FILLER_6_222 ();
 sg13g2_decap_4 FILLER_6_237 ();
 sg13g2_decap_4 FILLER_6_281 ();
 sg13g2_decap_4 FILLER_6_295 ();
 sg13g2_fill_2 FILLER_6_314 ();
 sg13g2_decap_4 FILLER_6_326 ();
 sg13g2_fill_1 FILLER_6_360 ();
 sg13g2_fill_1 FILLER_6_390 ();
 sg13g2_fill_1 FILLER_6_395 ();
 sg13g2_fill_1 FILLER_7_0 ();
 sg13g2_decap_4 FILLER_7_47 ();
 sg13g2_decap_4 FILLER_7_98 ();
 sg13g2_fill_1 FILLER_7_115 ();
 sg13g2_fill_2 FILLER_7_126 ();
 sg13g2_decap_8 FILLER_7_203 ();
 sg13g2_fill_2 FILLER_7_210 ();
 sg13g2_fill_1 FILLER_7_212 ();
 sg13g2_decap_8 FILLER_7_227 ();
 sg13g2_fill_2 FILLER_7_279 ();
 sg13g2_fill_2 FILLER_7_331 ();
 sg13g2_fill_1 FILLER_7_333 ();
 sg13g2_fill_2 FILLER_7_374 ();
 sg13g2_fill_1 FILLER_7_376 ();
 sg13g2_fill_2 FILLER_8_0 ();
 sg13g2_fill_1 FILLER_8_2 ();
 sg13g2_fill_2 FILLER_8_20 ();
 sg13g2_fill_1 FILLER_8_60 ();
 sg13g2_fill_2 FILLER_8_71 ();
 sg13g2_fill_2 FILLER_8_97 ();
 sg13g2_fill_2 FILLER_8_149 ();
 sg13g2_fill_1 FILLER_8_151 ();
 sg13g2_fill_2 FILLER_8_157 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_fill_2 FILLER_8_180 ();
 sg13g2_decap_4 FILLER_8_202 ();
 sg13g2_fill_1 FILLER_8_206 ();
 sg13g2_decap_8 FILLER_8_227 ();
 sg13g2_decap_8 FILLER_8_234 ();
 sg13g2_fill_2 FILLER_8_241 ();
 sg13g2_fill_1 FILLER_8_253 ();
 sg13g2_fill_2 FILLER_8_259 ();
 sg13g2_fill_1 FILLER_8_261 ();
 sg13g2_fill_2 FILLER_8_267 ();
 sg13g2_fill_2 FILLER_8_304 ();
 sg13g2_fill_1 FILLER_8_316 ();
 sg13g2_fill_2 FILLER_8_327 ();
 sg13g2_fill_2 FILLER_8_349 ();
 sg13g2_fill_1 FILLER_8_351 ();
 sg13g2_fill_1 FILLER_8_391 ();
 sg13g2_fill_2 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_72 ();
 sg13g2_decap_4 FILLER_9_102 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_194 ();
 sg13g2_decap_8 FILLER_9_201 ();
 sg13g2_decap_8 FILLER_9_208 ();
 sg13g2_fill_2 FILLER_9_229 ();
 sg13g2_fill_1 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_297 ();
 sg13g2_fill_2 FILLER_9_304 ();
 sg13g2_decap_8 FILLER_9_311 ();
 sg13g2_decap_4 FILLER_9_318 ();
 sg13g2_fill_1 FILLER_9_335 ();
 sg13g2_fill_2 FILLER_9_344 ();
 sg13g2_fill_1 FILLER_9_346 ();
 sg13g2_decap_8 FILLER_9_352 ();
 sg13g2_fill_1 FILLER_9_359 ();
 sg13g2_fill_1 FILLER_9_380 ();
 sg13g2_fill_2 FILLER_10_31 ();
 sg13g2_fill_2 FILLER_10_43 ();
 sg13g2_fill_2 FILLER_10_59 ();
 sg13g2_fill_1 FILLER_10_61 ();
 sg13g2_fill_2 FILLER_10_116 ();
 sg13g2_fill_1 FILLER_10_118 ();
 sg13g2_fill_2 FILLER_10_124 ();
 sg13g2_fill_1 FILLER_10_139 ();
 sg13g2_fill_2 FILLER_10_163 ();
 sg13g2_decap_4 FILLER_10_202 ();
 sg13g2_fill_2 FILLER_10_206 ();
 sg13g2_fill_1 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_233 ();
 sg13g2_fill_2 FILLER_10_240 ();
 sg13g2_fill_2 FILLER_10_252 ();
 sg13g2_fill_1 FILLER_10_259 ();
 sg13g2_fill_1 FILLER_10_280 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_fill_2 FILLER_10_321 ();
 sg13g2_fill_1 FILLER_11_0 ();
 sg13g2_fill_1 FILLER_11_9 ();
 sg13g2_fill_2 FILLER_11_14 ();
 sg13g2_fill_2 FILLER_11_66 ();
 sg13g2_fill_2 FILLER_11_113 ();
 sg13g2_fill_1 FILLER_11_130 ();
 sg13g2_fill_2 FILLER_11_154 ();
 sg13g2_fill_1 FILLER_11_156 ();
 sg13g2_fill_1 FILLER_11_162 ();
 sg13g2_fill_2 FILLER_11_173 ();
 sg13g2_fill_1 FILLER_11_175 ();
 sg13g2_decap_4 FILLER_11_210 ();
 sg13g2_decap_4 FILLER_11_299 ();
 sg13g2_decap_4 FILLER_11_335 ();
 sg13g2_fill_1 FILLER_11_339 ();
 sg13g2_decap_4 FILLER_11_345 ();
 sg13g2_fill_1 FILLER_11_349 ();
 sg13g2_fill_2 FILLER_11_355 ();
 sg13g2_fill_1 FILLER_11_357 ();
 sg13g2_fill_1 FILLER_11_367 ();
 sg13g2_fill_1 FILLER_11_378 ();
 sg13g2_fill_2 FILLER_11_389 ();
 sg13g2_fill_1 FILLER_11_391 ();
 sg13g2_fill_1 FILLER_12_0 ();
 sg13g2_fill_2 FILLER_12_19 ();
 sg13g2_fill_1 FILLER_12_21 ();
 sg13g2_fill_1 FILLER_12_58 ();
 sg13g2_fill_2 FILLER_12_91 ();
 sg13g2_fill_1 FILLER_12_93 ();
 sg13g2_fill_2 FILLER_12_171 ();
 sg13g2_fill_2 FILLER_12_177 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_205 ();
 sg13g2_fill_1 FILLER_12_207 ();
 sg13g2_decap_4 FILLER_12_223 ();
 sg13g2_fill_1 FILLER_12_227 ();
 sg13g2_fill_2 FILLER_12_233 ();
 sg13g2_fill_1 FILLER_12_235 ();
 sg13g2_fill_2 FILLER_12_240 ();
 sg13g2_fill_1 FILLER_12_242 ();
 sg13g2_fill_1 FILLER_12_248 ();
 sg13g2_fill_2 FILLER_12_264 ();
 sg13g2_decap_8 FILLER_12_286 ();
 sg13g2_decap_8 FILLER_12_293 ();
 sg13g2_fill_2 FILLER_12_300 ();
 sg13g2_fill_2 FILLER_12_312 ();
 sg13g2_fill_1 FILLER_12_314 ();
 sg13g2_fill_1 FILLER_12_318 ();
 sg13g2_decap_4 FILLER_12_329 ();
 sg13g2_fill_1 FILLER_12_348 ();
 sg13g2_fill_2 FILLER_12_379 ();
 sg13g2_fill_1 FILLER_12_381 ();
 sg13g2_fill_2 FILLER_13_0 ();
 sg13g2_fill_2 FILLER_13_103 ();
 sg13g2_fill_1 FILLER_13_105 ();
 sg13g2_fill_2 FILLER_13_121 ();
 sg13g2_fill_2 FILLER_13_181 ();
 sg13g2_fill_1 FILLER_13_183 ();
 sg13g2_decap_4 FILLER_13_197 ();
 sg13g2_fill_2 FILLER_13_219 ();
 sg13g2_fill_1 FILLER_13_221 ();
 sg13g2_decap_4 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_291 ();
 sg13g2_fill_2 FILLER_13_372 ();
 sg13g2_fill_1 FILLER_13_408 ();
 sg13g2_fill_1 FILLER_14_0 ();
 sg13g2_fill_2 FILLER_14_47 ();
 sg13g2_fill_1 FILLER_14_93 ();
 sg13g2_fill_2 FILLER_14_99 ();
 sg13g2_fill_2 FILLER_14_115 ();
 sg13g2_fill_1 FILLER_14_151 ();
 sg13g2_fill_1 FILLER_14_184 ();
 sg13g2_decap_4 FILLER_14_190 ();
 sg13g2_fill_2 FILLER_14_194 ();
 sg13g2_fill_2 FILLER_14_216 ();
 sg13g2_decap_8 FILLER_14_230 ();
 sg13g2_decap_8 FILLER_14_237 ();
 sg13g2_decap_4 FILLER_14_244 ();
 sg13g2_fill_2 FILLER_14_253 ();
 sg13g2_decap_4 FILLER_14_260 ();
 sg13g2_fill_1 FILLER_14_264 ();
 sg13g2_decap_8 FILLER_14_285 ();
 sg13g2_fill_2 FILLER_14_292 ();
 sg13g2_decap_4 FILLER_14_306 ();
 sg13g2_decap_4 FILLER_14_323 ();
 sg13g2_fill_2 FILLER_14_332 ();
 sg13g2_fill_1 FILLER_14_334 ();
 sg13g2_fill_2 FILLER_14_339 ();
 sg13g2_decap_8 FILLER_14_346 ();
 sg13g2_fill_2 FILLER_14_353 ();
 sg13g2_fill_1 FILLER_14_355 ();
 sg13g2_fill_2 FILLER_14_366 ();
 sg13g2_fill_2 FILLER_14_378 ();
 sg13g2_fill_1 FILLER_14_380 ();
 sg13g2_fill_2 FILLER_15_32 ();
 sg13g2_fill_1 FILLER_15_34 ();
 sg13g2_fill_2 FILLER_15_55 ();
 sg13g2_fill_2 FILLER_15_107 ();
 sg13g2_fill_2 FILLER_15_188 ();
 sg13g2_fill_1 FILLER_15_190 ();
 sg13g2_fill_2 FILLER_15_195 ();
 sg13g2_fill_2 FILLER_15_206 ();
 sg13g2_decap_8 FILLER_15_213 ();
 sg13g2_decap_8 FILLER_15_220 ();
 sg13g2_fill_1 FILLER_15_227 ();
 sg13g2_fill_2 FILLER_15_233 ();
 sg13g2_fill_1 FILLER_15_235 ();
 sg13g2_fill_1 FILLER_15_286 ();
 sg13g2_fill_2 FILLER_15_313 ();
 sg13g2_fill_1 FILLER_15_315 ();
 sg13g2_fill_2 FILLER_15_407 ();
 sg13g2_fill_2 FILLER_16_0 ();
 sg13g2_fill_1 FILLER_16_2 ();
 sg13g2_fill_1 FILLER_16_20 ();
 sg13g2_fill_2 FILLER_16_25 ();
 sg13g2_fill_1 FILLER_16_27 ();
 sg13g2_fill_2 FILLER_16_44 ();
 sg13g2_fill_2 FILLER_16_84 ();
 sg13g2_fill_1 FILLER_16_86 ();
 sg13g2_fill_1 FILLER_16_124 ();
 sg13g2_fill_2 FILLER_16_156 ();
 sg13g2_fill_1 FILLER_16_158 ();
 sg13g2_fill_2 FILLER_16_199 ();
 sg13g2_fill_1 FILLER_16_206 ();
 sg13g2_decap_8 FILLER_16_241 ();
 sg13g2_fill_2 FILLER_16_248 ();
 sg13g2_decap_4 FILLER_16_260 ();
 sg13g2_fill_2 FILLER_16_264 ();
 sg13g2_fill_2 FILLER_16_271 ();
 sg13g2_fill_1 FILLER_16_293 ();
 sg13g2_decap_8 FILLER_16_321 ();
 sg13g2_fill_1 FILLER_16_328 ();
 sg13g2_decap_8 FILLER_16_334 ();
 sg13g2_fill_1 FILLER_16_341 ();
 sg13g2_fill_2 FILLER_16_347 ();
 sg13g2_fill_1 FILLER_16_359 ();
 sg13g2_fill_1 FILLER_16_380 ();
 sg13g2_fill_2 FILLER_17_0 ();
 sg13g2_fill_1 FILLER_17_2 ();
 sg13g2_fill_2 FILLER_17_34 ();
 sg13g2_fill_1 FILLER_17_36 ();
 sg13g2_fill_2 FILLER_17_61 ();
 sg13g2_fill_1 FILLER_17_97 ();
 sg13g2_fill_2 FILLER_17_104 ();
 sg13g2_fill_1 FILLER_17_106 ();
 sg13g2_fill_2 FILLER_17_153 ();
 sg13g2_fill_2 FILLER_17_173 ();
 sg13g2_fill_1 FILLER_17_192 ();
 sg13g2_fill_1 FILLER_17_202 ();
 sg13g2_decap_8 FILLER_17_210 ();
 sg13g2_decap_8 FILLER_17_217 ();
 sg13g2_fill_2 FILLER_17_224 ();
 sg13g2_decap_8 FILLER_17_236 ();
 sg13g2_fill_1 FILLER_17_253 ();
 sg13g2_decap_4 FILLER_17_259 ();
 sg13g2_decap_4 FILLER_17_273 ();
 sg13g2_fill_2 FILLER_17_277 ();
 sg13g2_decap_4 FILLER_17_284 ();
 sg13g2_fill_2 FILLER_17_288 ();
 sg13g2_fill_1 FILLER_17_305 ();
 sg13g2_decap_4 FILLER_17_318 ();
 sg13g2_fill_2 FILLER_17_387 ();
 sg13g2_fill_1 FILLER_17_389 ();
 sg13g2_fill_2 FILLER_17_406 ();
 sg13g2_fill_1 FILLER_17_408 ();
 sg13g2_fill_2 FILLER_18_0 ();
 sg13g2_fill_1 FILLER_18_2 ();
 sg13g2_fill_2 FILLER_18_60 ();
 sg13g2_fill_1 FILLER_18_77 ();
 sg13g2_fill_2 FILLER_18_110 ();
 sg13g2_fill_1 FILLER_18_112 ();
 sg13g2_fill_1 FILLER_18_124 ();
 sg13g2_fill_1 FILLER_18_145 ();
 sg13g2_fill_2 FILLER_18_150 ();
 sg13g2_fill_1 FILLER_18_152 ();
 sg13g2_fill_2 FILLER_18_170 ();
 sg13g2_fill_1 FILLER_18_172 ();
 sg13g2_fill_2 FILLER_18_179 ();
 sg13g2_fill_1 FILLER_18_191 ();
 sg13g2_fill_1 FILLER_18_200 ();
 sg13g2_fill_1 FILLER_18_205 ();
 sg13g2_decap_8 FILLER_18_216 ();
 sg13g2_fill_1 FILLER_18_238 ();
 sg13g2_fill_2 FILLER_18_319 ();
 sg13g2_fill_1 FILLER_18_364 ();
 sg13g2_fill_1 FILLER_18_380 ();
 sg13g2_fill_1 FILLER_19_126 ();
 sg13g2_fill_1 FILLER_19_136 ();
 sg13g2_fill_2 FILLER_19_145 ();
 sg13g2_fill_2 FILLER_19_175 ();
 sg13g2_fill_1 FILLER_19_181 ();
 sg13g2_fill_2 FILLER_19_201 ();
 sg13g2_fill_2 FILLER_19_212 ();
 sg13g2_fill_2 FILLER_19_218 ();
 sg13g2_fill_2 FILLER_19_250 ();
 sg13g2_fill_1 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_fill_1 FILLER_19_280 ();
 sg13g2_decap_4 FILLER_19_286 ();
 sg13g2_fill_2 FILLER_19_307 ();
 sg13g2_decap_4 FILLER_19_317 ();
 sg13g2_fill_2 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_328 ();
 sg13g2_fill_2 FILLER_19_338 ();
 sg13g2_fill_2 FILLER_19_372 ();
 sg13g2_fill_1 FILLER_20_0 ();
 sg13g2_fill_2 FILLER_20_17 ();
 sg13g2_fill_1 FILLER_20_19 ();
 sg13g2_fill_2 FILLER_20_39 ();
 sg13g2_fill_1 FILLER_20_41 ();
 sg13g2_fill_2 FILLER_20_88 ();
 sg13g2_fill_1 FILLER_20_90 ();
 sg13g2_fill_2 FILLER_20_174 ();
 sg13g2_fill_1 FILLER_20_176 ();
 sg13g2_fill_2 FILLER_20_189 ();
 sg13g2_decap_8 FILLER_20_234 ();
 sg13g2_decap_4 FILLER_20_241 ();
 sg13g2_fill_1 FILLER_20_368 ();
 sg13g2_fill_2 FILLER_21_0 ();
 sg13g2_fill_1 FILLER_21_2 ();
 sg13g2_fill_1 FILLER_21_48 ();
 sg13g2_fill_1 FILLER_21_103 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_fill_2 FILLER_21_177 ();
 sg13g2_decap_4 FILLER_21_242 ();
 sg13g2_fill_1 FILLER_21_262 ();
 sg13g2_fill_1 FILLER_21_285 ();
 sg13g2_decap_4 FILLER_21_291 ();
 sg13g2_fill_1 FILLER_21_300 ();
 sg13g2_fill_2 FILLER_21_305 ();
 sg13g2_fill_1 FILLER_21_307 ();
 sg13g2_fill_1 FILLER_21_362 ();
 sg13g2_fill_2 FILLER_21_373 ();
 sg13g2_fill_2 FILLER_21_384 ();
 sg13g2_fill_1 FILLER_21_386 ();
 sg13g2_fill_1 FILLER_21_391 ();
 sg13g2_fill_1 FILLER_22_0 ();
 sg13g2_fill_2 FILLER_22_19 ();
 sg13g2_fill_1 FILLER_22_43 ();
 sg13g2_fill_2 FILLER_22_58 ();
 sg13g2_fill_1 FILLER_22_93 ();
 sg13g2_fill_2 FILLER_22_107 ();
 sg13g2_fill_1 FILLER_22_109 ();
 sg13g2_fill_1 FILLER_22_156 ();
 sg13g2_fill_1 FILLER_22_171 ();
 sg13g2_fill_1 FILLER_22_189 ();
 sg13g2_fill_2 FILLER_22_210 ();
 sg13g2_fill_1 FILLER_22_246 ();
 sg13g2_fill_2 FILLER_22_260 ();
 sg13g2_fill_1 FILLER_22_275 ();
 sg13g2_fill_1 FILLER_22_289 ();
 sg13g2_decap_4 FILLER_22_294 ();
 sg13g2_fill_1 FILLER_22_298 ();
 sg13g2_fill_1 FILLER_22_329 ();
 sg13g2_fill_1 FILLER_22_353 ();
 sg13g2_fill_2 FILLER_22_366 ();
 sg13g2_fill_1 FILLER_22_368 ();
 sg13g2_fill_1 FILLER_23_0 ();
 sg13g2_fill_2 FILLER_23_62 ();
 sg13g2_fill_1 FILLER_23_64 ();
 sg13g2_fill_2 FILLER_23_73 ();
 sg13g2_fill_1 FILLER_23_75 ();
 sg13g2_fill_1 FILLER_23_81 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_183 ();
 sg13g2_fill_1 FILLER_23_189 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_2 FILLER_23_247 ();
 sg13g2_fill_1 FILLER_23_271 ();
 sg13g2_decap_4 FILLER_23_277 ();
 sg13g2_fill_1 FILLER_23_281 ();
 sg13g2_fill_2 FILLER_23_382 ();
 sg13g2_fill_2 FILLER_23_407 ();
 sg13g2_fill_2 FILLER_24_88 ();
 sg13g2_fill_1 FILLER_24_90 ();
 sg13g2_fill_2 FILLER_24_103 ();
 sg13g2_fill_2 FILLER_24_129 ();
 sg13g2_fill_2 FILLER_24_175 ();
 sg13g2_fill_1 FILLER_24_188 ();
 sg13g2_fill_2 FILLER_24_200 ();
 sg13g2_fill_1 FILLER_24_213 ();
 sg13g2_fill_1 FILLER_24_242 ();
 sg13g2_fill_1 FILLER_24_264 ();
 sg13g2_fill_2 FILLER_24_278 ();
 sg13g2_fill_1 FILLER_24_318 ();
 sg13g2_fill_2 FILLER_24_331 ();
 sg13g2_fill_1 FILLER_24_333 ();
 sg13g2_fill_1 FILLER_24_349 ();
 sg13g2_fill_1 FILLER_25_0 ();
 sg13g2_fill_2 FILLER_25_86 ();
 sg13g2_fill_1 FILLER_25_101 ();
 sg13g2_fill_2 FILLER_25_113 ();
 sg13g2_fill_1 FILLER_25_115 ();
 sg13g2_fill_1 FILLER_25_132 ();
 sg13g2_fill_2 FILLER_25_138 ();
 sg13g2_fill_1 FILLER_25_140 ();
 sg13g2_fill_2 FILLER_25_185 ();
 sg13g2_fill_2 FILLER_25_200 ();
 sg13g2_fill_1 FILLER_25_202 ();
 sg13g2_fill_2 FILLER_25_225 ();
 sg13g2_fill_1 FILLER_25_248 ();
 sg13g2_fill_2 FILLER_25_260 ();
 sg13g2_fill_2 FILLER_25_278 ();
 sg13g2_fill_1 FILLER_25_280 ();
 sg13g2_fill_2 FILLER_25_334 ();
 sg13g2_fill_2 FILLER_25_386 ();
 sg13g2_fill_1 FILLER_25_401 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_fill_1 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_56 ();
 sg13g2_fill_2 FILLER_26_78 ();
 sg13g2_fill_1 FILLER_26_80 ();
 sg13g2_fill_1 FILLER_26_99 ();
 sg13g2_fill_2 FILLER_26_118 ();
 sg13g2_fill_1 FILLER_26_150 ();
 sg13g2_fill_2 FILLER_26_156 ();
 sg13g2_fill_1 FILLER_26_158 ();
 sg13g2_fill_1 FILLER_26_211 ();
 sg13g2_fill_1 FILLER_26_244 ();
 sg13g2_fill_1 FILLER_26_250 ();
 sg13g2_fill_2 FILLER_26_261 ();
 sg13g2_fill_2 FILLER_26_274 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_fill_2 FILLER_26_297 ();
 sg13g2_fill_1 FILLER_26_317 ();
 sg13g2_fill_2 FILLER_27_29 ();
 sg13g2_fill_2 FILLER_27_49 ();
 sg13g2_fill_1 FILLER_27_51 ();
 sg13g2_fill_2 FILLER_27_68 ();
 sg13g2_fill_2 FILLER_27_76 ();
 sg13g2_fill_1 FILLER_27_103 ();
 sg13g2_fill_1 FILLER_27_153 ();
 sg13g2_fill_2 FILLER_27_248 ();
 sg13g2_fill_1 FILLER_27_390 ();
 sg13g2_fill_2 FILLER_28_61 ();
 sg13g2_fill_1 FILLER_28_63 ();
 sg13g2_fill_2 FILLER_28_114 ();
 sg13g2_fill_1 FILLER_28_116 ();
 sg13g2_fill_2 FILLER_28_156 ();
 sg13g2_fill_1 FILLER_28_158 ();
 sg13g2_fill_2 FILLER_28_178 ();
 sg13g2_fill_2 FILLER_28_200 ();
 sg13g2_fill_1 FILLER_28_202 ();
 sg13g2_fill_2 FILLER_28_221 ();
 sg13g2_fill_1 FILLER_28_223 ();
 sg13g2_fill_2 FILLER_28_242 ();
 sg13g2_fill_2 FILLER_28_249 ();
 sg13g2_fill_2 FILLER_28_279 ();
 sg13g2_fill_1 FILLER_28_281 ();
 sg13g2_fill_1 FILLER_28_297 ();
 sg13g2_fill_1 FILLER_28_336 ();
 sg13g2_fill_1 FILLER_28_355 ();
 sg13g2_fill_1 FILLER_29_50 ();
 sg13g2_fill_2 FILLER_29_83 ();
 sg13g2_fill_2 FILLER_29_111 ();
 sg13g2_fill_2 FILLER_29_134 ();
 sg13g2_fill_1 FILLER_29_136 ();
 sg13g2_fill_2 FILLER_29_142 ();
 sg13g2_fill_1 FILLER_29_155 ();
 sg13g2_fill_2 FILLER_29_248 ();
 sg13g2_fill_1 FILLER_29_250 ();
 sg13g2_fill_2 FILLER_29_274 ();
 sg13g2_fill_1 FILLER_29_276 ();
 sg13g2_fill_1 FILLER_29_296 ();
 sg13g2_fill_1 FILLER_29_319 ();
 sg13g2_fill_2 FILLER_29_325 ();
 sg13g2_fill_2 FILLER_29_407 ();
 sg13g2_fill_1 FILLER_30_0 ();
 sg13g2_fill_2 FILLER_30_75 ();
 sg13g2_fill_1 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_126 ();
 sg13g2_fill_1 FILLER_30_237 ();
 sg13g2_fill_2 FILLER_30_251 ();
 sg13g2_fill_1 FILLER_30_253 ();
 sg13g2_fill_2 FILLER_30_279 ();
 sg13g2_fill_1 FILLER_30_281 ();
 sg13g2_fill_1 FILLER_30_301 ();
 sg13g2_fill_1 FILLER_30_375 ();
 sg13g2_fill_1 FILLER_31_72 ();
 sg13g2_fill_2 FILLER_31_78 ();
 sg13g2_fill_1 FILLER_31_103 ();
 sg13g2_fill_2 FILLER_31_135 ();
 sg13g2_fill_1 FILLER_31_137 ();
 sg13g2_fill_1 FILLER_31_160 ();
 sg13g2_fill_1 FILLER_31_253 ();
 sg13g2_fill_2 FILLER_31_283 ();
 sg13g2_fill_2 FILLER_31_290 ();
 sg13g2_fill_1 FILLER_31_292 ();
 sg13g2_fill_1 FILLER_31_298 ();
 sg13g2_fill_2 FILLER_31_332 ();
 sg13g2_fill_2 FILLER_31_344 ();
 sg13g2_fill_2 FILLER_31_351 ();
 sg13g2_fill_2 FILLER_31_376 ();
 sg13g2_fill_2 FILLER_32_37 ();
 sg13g2_fill_1 FILLER_32_39 ();
 sg13g2_fill_2 FILLER_32_104 ();
 sg13g2_fill_2 FILLER_32_119 ();
 sg13g2_fill_1 FILLER_32_121 ();
 sg13g2_fill_2 FILLER_32_135 ();
 sg13g2_fill_1 FILLER_32_137 ();
 sg13g2_fill_2 FILLER_32_171 ();
 sg13g2_fill_1 FILLER_32_191 ();
 sg13g2_fill_2 FILLER_32_202 ();
 sg13g2_fill_1 FILLER_32_204 ();
 sg13g2_fill_1 FILLER_32_232 ();
 sg13g2_fill_1 FILLER_32_243 ();
 sg13g2_fill_2 FILLER_32_290 ();
 sg13g2_fill_1 FILLER_32_322 ();
 sg13g2_fill_2 FILLER_32_406 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_1 FILLER_33_0 ();
 sg13g2_fill_2 FILLER_33_29 ();
 sg13g2_fill_2 FILLER_33_59 ();
 sg13g2_fill_1 FILLER_33_61 ();
 sg13g2_fill_1 FILLER_33_95 ();
 sg13g2_fill_2 FILLER_33_127 ();
 sg13g2_fill_1 FILLER_33_129 ();
 sg13g2_fill_1 FILLER_33_139 ();
 sg13g2_fill_1 FILLER_33_160 ();
 sg13g2_fill_2 FILLER_33_232 ();
 sg13g2_fill_1 FILLER_33_244 ();
 sg13g2_fill_1 FILLER_34_23 ();
 sg13g2_fill_2 FILLER_34_47 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_fill_2 FILLER_34_59 ();
 sg13g2_fill_1 FILLER_34_71 ();
 sg13g2_fill_1 FILLER_34_101 ();
 sg13g2_fill_2 FILLER_34_142 ();
 sg13g2_fill_2 FILLER_34_194 ();
 sg13g2_fill_1 FILLER_34_196 ();
 sg13g2_fill_2 FILLER_34_207 ();
 sg13g2_fill_1 FILLER_34_209 ();
 sg13g2_fill_2 FILLER_34_253 ();
 sg13g2_fill_2 FILLER_34_273 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_fill_2 FILLER_34_311 ();
 sg13g2_fill_1 FILLER_34_313 ();
 sg13g2_fill_1 FILLER_34_344 ();
 sg13g2_fill_2 FILLER_34_360 ();
 sg13g2_fill_1 FILLER_34_380 ();
 sg13g2_fill_2 FILLER_35_263 ();
 sg13g2_fill_1 FILLER_35_265 ();
 sg13g2_fill_2 FILLER_35_306 ();
 sg13g2_fill_1 FILLER_35_318 ();
 sg13g2_fill_2 FILLER_36_0 ();
 sg13g2_fill_1 FILLER_36_2 ();
 sg13g2_fill_1 FILLER_36_64 ();
 sg13g2_fill_1 FILLER_36_89 ();
 sg13g2_fill_2 FILLER_36_152 ();
 sg13g2_fill_2 FILLER_36_222 ();
 sg13g2_fill_1 FILLER_36_248 ();
 sg13g2_fill_1 FILLER_36_332 ();
 sg13g2_fill_1 FILLER_36_346 ();
 sg13g2_fill_2 FILLER_37_0 ();
 sg13g2_fill_1 FILLER_37_2 ();
 sg13g2_fill_2 FILLER_37_49 ();
 sg13g2_fill_1 FILLER_37_51 ();
 sg13g2_fill_2 FILLER_37_127 ();
 sg13g2_fill_1 FILLER_37_129 ();
 sg13g2_fill_2 FILLER_37_139 ();
 sg13g2_fill_2 FILLER_37_212 ();
 sg13g2_fill_2 FILLER_37_260 ();
 sg13g2_fill_1 FILLER_37_262 ();
 sg13g2_fill_1 FILLER_37_277 ();
 sg13g2_fill_2 FILLER_37_394 ();
 sg13g2_fill_1 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_54 ();
 sg13g2_fill_2 FILLER_38_70 ();
 sg13g2_fill_2 FILLER_38_281 ();
 sg13g2_fill_1 FILLER_38_283 ();
 sg13g2_fill_1 FILLER_38_338 ();
 sg13g2_fill_2 FILLER_38_376 ();
endmodule
