module tt_um_rebeccargb_vga_pride (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire clknet_0_clk;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \flag.flag_abrosexual_inst.pix_x[0] ;
 wire \flag.flag_abrosexual_inst.pix_x[1] ;
 wire \flag.flag_abrosexual_inst.pix_x[2] ;
 wire \flag.flag_abrosexual_inst.pix_x[3] ;
 wire \flag.flag_abrosexual_inst.pix_x[4] ;
 wire \flag.flag_abrosexual_inst.pix_x[5] ;
 wire \flag.flag_abrosexual_inst.pix_x[6] ;
 wire \flag.flag_abrosexual_inst.pix_x[7] ;
 wire \flag.flag_abrosexual_inst.pix_x[8] ;
 wire \flag.flag_abrosexual_inst.pix_x[9] ;
 wire \flag.flag_abrosexual_inst.pix_y[0] ;
 wire \flag.flag_abrosexual_inst.pix_y[1] ;
 wire \flag.flag_abrosexual_inst.pix_y[2] ;
 wire \flag.flag_abrosexual_inst.pix_y[3] ;
 wire \flag.flag_abrosexual_inst.pix_y[4] ;
 wire \flag.flag_abrosexual_inst.pix_y[5] ;
 wire \flag.flag_abrosexual_inst.pix_y[6] ;
 wire \flag.flag_abrosexual_inst.pix_y[7] ;
 wire \flag.flag_abrosexual_inst.pix_y[8] ;
 wire hsync;
 wire \hvsync_gen.vpos[9] ;
 wire \hvsync_gen.vsync ;
 wire \reset_latch[0] ;
 wire \reset_latch[1] ;
 wire \reset_latch[2] ;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;

 sg13g2_inv_1 _2778_ (.Y(_2558_),
    .A(net569));
 sg13g2_inv_4 _2779_ (.A(net575),
    .Y(_2569_));
 sg13g2_inv_4 _2780_ (.A(net584),
    .Y(_2580_));
 sg13g2_inv_4 _2781_ (.A(net587),
    .Y(_2591_));
 sg13g2_inv_1 _2782_ (.Y(_2602_),
    .A(net593));
 sg13g2_inv_8 _2783_ (.Y(_2613_),
    .A(net595));
 sg13g2_inv_4 _2784_ (.A(net598),
    .Y(_2624_));
 sg13g2_inv_8 _2785_ (.Y(_2635_),
    .A(net602));
 sg13g2_inv_2 _2786_ (.Y(_2646_),
    .A(net653));
 sg13g2_inv_1 _2787_ (.Y(_2657_),
    .A(net4));
 sg13g2_inv_2 _2788_ (.Y(_2668_),
    .A(net645));
 sg13g2_inv_2 _2789_ (.Y(_2679_),
    .A(net636));
 sg13g2_inv_4 _2790_ (.A(net641),
    .Y(_2690_));
 sg13g2_inv_2 _2791_ (.Y(_2701_),
    .A(net632));
 sg13g2_inv_4 _2792_ (.A(net623),
    .Y(_2712_));
 sg13g2_inv_1 _2793_ (.Y(_2723_),
    .A(net617));
 sg13g2_inv_1 _2794_ (.Y(_2734_),
    .A(net613));
 sg13g2_inv_2 _2795_ (.Y(_2745_),
    .A(net608));
 sg13g2_inv_1 _2796_ (.Y(_0032_),
    .A(\reset_latch[2] ));
 sg13g2_inv_4 _2797_ (.A(net656),
    .Y(_0043_));
 sg13g2_inv_2 _2798_ (.Y(_0054_),
    .A(\counter[3] ));
 sg13g2_mux2_1 _2799_ (.A0(\counter[6] ),
    .A1(net12),
    .S(net1),
    .X(_0065_));
 sg13g2_mux2_1 _2800_ (.A0(\counter[5] ),
    .A1(net11),
    .S(net1),
    .X(_0076_));
 sg13g2_mux2_1 _2801_ (.A0(\counter[4] ),
    .A1(net10),
    .S(net1),
    .X(_0087_));
 sg13g2_nor2b_2 _2802_ (.A(_0076_),
    .B_N(_0087_),
    .Y(_0098_));
 sg13g2_nand2_2 _2803_ (.Y(_0109_),
    .A(net550),
    .B(_0098_));
 sg13g2_nand2_1 _2804_ (.Y(_0120_),
    .A(net9),
    .B(net1));
 sg13g2_o21ai_1 _2805_ (.B1(_0120_),
    .Y(_0131_),
    .A1(_0054_),
    .A2(net1));
 sg13g2_mux2_1 _2806_ (.A0(\counter[2] ),
    .A1(net8),
    .S(net1),
    .X(_0142_));
 sg13g2_nor2_2 _2807_ (.A(_0131_),
    .B(_0142_),
    .Y(_0153_));
 sg13g2_or2_1 _2808_ (.X(_0164_),
    .B(_0142_),
    .A(_0131_));
 sg13g2_mux2_1 _2809_ (.A0(\counter[1] ),
    .A1(net7),
    .S(net1),
    .X(_0175_));
 sg13g2_inv_1 _2810_ (.Y(_0186_),
    .A(_0175_));
 sg13g2_mux2_1 _2811_ (.A0(\counter[0] ),
    .A1(net6),
    .S(net1),
    .X(_0197_));
 sg13g2_nor2b_2 _2812_ (.A(_0175_),
    .B_N(_0197_),
    .Y(_0208_));
 sg13g2_and2_1 _2813_ (.A(_0153_),
    .B(_0208_),
    .X(_0219_));
 sg13g2_nand2_1 _2814_ (.Y(_0230_),
    .A(_0153_),
    .B(_0208_));
 sg13g2_nand2b_1 _2815_ (.Y(_0241_),
    .B(_0219_),
    .A_N(net516));
 sg13g2_nor2_2 _2816_ (.A(_0175_),
    .B(_0197_),
    .Y(_0252_));
 sg13g2_nor2b_2 _2817_ (.A(_0131_),
    .B_N(_0142_),
    .Y(_0263_));
 sg13g2_nand2_2 _2818_ (.Y(_0274_),
    .A(_0252_),
    .B(_0263_));
 sg13g2_nor2_2 _2819_ (.A(net516),
    .B(_0274_),
    .Y(_0285_));
 sg13g2_and2_1 _2820_ (.A(_0175_),
    .B(_0197_),
    .X(_0296_));
 sg13g2_nand2_2 _2821_ (.Y(_0307_),
    .A(_0153_),
    .B(_0296_));
 sg13g2_nor2_2 _2822_ (.A(net516),
    .B(_0307_),
    .Y(_0318_));
 sg13g2_or2_1 _2823_ (.X(_0329_),
    .B(_0307_),
    .A(net516));
 sg13g2_nand2_2 _2824_ (.Y(_0340_),
    .A(_0153_),
    .B(_0252_));
 sg13g2_nor2_2 _2825_ (.A(net516),
    .B(_0340_),
    .Y(_0351_));
 sg13g2_and2_1 _2826_ (.A(_0208_),
    .B(_0263_),
    .X(_0362_));
 sg13g2_nand2_2 _2827_ (.Y(_0373_),
    .A(_0208_),
    .B(_0263_));
 sg13g2_nor2_1 _2828_ (.A(net516),
    .B(_0373_),
    .Y(_0384_));
 sg13g2_nand2b_1 _2829_ (.Y(_0395_),
    .B(_0362_),
    .A_N(net516));
 sg13g2_nor2_2 _2830_ (.A(_0351_),
    .B(_0384_),
    .Y(_0406_));
 sg13g2_nor2_1 _2831_ (.A(_0076_),
    .B(_0087_),
    .Y(_0417_));
 sg13g2_inv_1 _2832_ (.Y(_0428_),
    .A(_0417_));
 sg13g2_nor2_2 _2833_ (.A(_0186_),
    .B(_0197_),
    .Y(_0439_));
 sg13g2_nand2_2 _2834_ (.Y(_0450_),
    .A(_0153_),
    .B(_0439_));
 sg13g2_nor2_2 _2835_ (.A(_0109_),
    .B(_0450_),
    .Y(_0461_));
 sg13g2_nand4_1 _2836_ (.B(_0241_),
    .C(_0406_),
    .A(net550),
    .Y(_0472_),
    .D(_0428_));
 sg13g2_nor4_1 _2837_ (.A(_0285_),
    .B(_0318_),
    .C(_0461_),
    .D(_0472_),
    .Y(_0483_));
 sg13g2_and2_1 _2838_ (.A(net573),
    .B(net577),
    .X(_0494_));
 sg13g2_nand2_1 _2839_ (.Y(_0505_),
    .A(net573),
    .B(net577));
 sg13g2_and2_1 _2840_ (.A(net577),
    .B(net583),
    .X(_0516_));
 sg13g2_nand2_2 _2841_ (.Y(_0527_),
    .A(net581),
    .B(net586));
 sg13g2_and3_1 _2842_ (.X(_0538_),
    .A(net573),
    .B(net578),
    .C(net582));
 sg13g2_nand3_1 _2843_ (.B(net580),
    .C(net586),
    .A(net576),
    .Y(_0549_));
 sg13g2_nor2_2 _2844_ (.A(net563),
    .B(_2569_),
    .Y(_0560_));
 sg13g2_nand2_1 _2845_ (.Y(_0571_),
    .A(net570),
    .B(net575));
 sg13g2_nor2_2 _2846_ (.A(_0527_),
    .B(net548),
    .Y(_0582_));
 sg13g2_inv_2 _2847_ (.Y(_0593_),
    .A(_0582_));
 sg13g2_nor2_2 _2848_ (.A(net618),
    .B(net612),
    .Y(_0604_));
 sg13g2_nand2_1 _2849_ (.Y(_0615_),
    .A(net554),
    .B(net552));
 sg13g2_nor2_1 _2850_ (.A(net551),
    .B(_0604_),
    .Y(_0626_));
 sg13g2_or4_1 _2851_ (.A(\hvsync_gen.vpos[9] ),
    .B(_0483_),
    .C(_0582_),
    .D(_0626_),
    .X(_0637_));
 sg13g2_nor2_2 _2852_ (.A(net622),
    .B(net616),
    .Y(_0648_));
 sg13g2_or2_1 _2853_ (.X(_0659_),
    .B(net617),
    .A(net623));
 sg13g2_o21ai_1 _2854_ (.B1(net611),
    .Y(_0670_),
    .A1(net623),
    .A2(net617));
 sg13g2_and2_1 _2855_ (.A(_2745_),
    .B(_0670_),
    .X(_0681_));
 sg13g2_nor2_1 _2856_ (.A(net643),
    .B(net639),
    .Y(_0692_));
 sg13g2_or2_1 _2857_ (.X(_0703_),
    .B(net645),
    .A(net650));
 sg13g2_nor3_2 _2858_ (.A(net652),
    .B(net646),
    .C(net642),
    .Y(_0714_));
 sg13g2_or3_1 _2859_ (.A(net652),
    .B(net646),
    .C(net642),
    .X(_0725_));
 sg13g2_nor2_2 _2860_ (.A(net638),
    .B(net641),
    .Y(_0736_));
 sg13g2_nand2_1 _2861_ (.Y(_0747_),
    .A(net558),
    .B(_2690_));
 sg13g2_or4_1 _2862_ (.A(net652),
    .B(\flag.flag_abrosexual_inst.pix_x[1] ),
    .C(net637),
    .D(net642),
    .X(_0758_));
 sg13g2_nand3_1 _2863_ (.B(_0670_),
    .C(_0758_),
    .A(net551),
    .Y(_0769_));
 sg13g2_xnor2_1 _2864_ (.Y(_0780_),
    .A(net634),
    .B(_0769_));
 sg13g2_xnor2_1 _2865_ (.Y(_0791_),
    .A(net557),
    .B(_0769_));
 sg13g2_nand3_1 _2866_ (.B(_0670_),
    .C(_0703_),
    .A(net551),
    .Y(_0802_));
 sg13g2_xnor2_1 _2867_ (.Y(_0813_),
    .A(_2690_),
    .B(_0802_));
 sg13g2_xnor2_1 _2868_ (.Y(_0824_),
    .A(net642),
    .B(_0802_));
 sg13g2_nor2_1 _2869_ (.A(net514),
    .B(net513),
    .Y(_0835_));
 sg13g2_nand2_1 _2870_ (.Y(_0846_),
    .A(net515),
    .B(net512));
 sg13g2_nand3_1 _2871_ (.B(_0670_),
    .C(_0725_),
    .A(net551),
    .Y(_0857_));
 sg13g2_xnor2_1 _2872_ (.Y(_0868_),
    .A(_2679_),
    .B(_0857_));
 sg13g2_xnor2_1 _2873_ (.Y(_0879_),
    .A(net638),
    .B(_0857_));
 sg13g2_a21oi_1 _2874_ (.A1(net513),
    .A2(net510),
    .Y(_0890_),
    .B1(_0835_));
 sg13g2_inv_1 _2875_ (.Y(_0901_),
    .A(_0890_));
 sg13g2_nor2_2 _2876_ (.A(net634),
    .B(net629),
    .Y(_0912_));
 sg13g2_or2_1 _2877_ (.X(_0923_),
    .B(net629),
    .A(net635));
 sg13g2_nor2_1 _2878_ (.A(net636),
    .B(net632),
    .Y(_0934_));
 sg13g2_or2_1 _2879_ (.X(_0945_),
    .B(net632),
    .A(net636));
 sg13g2_nor3_2 _2880_ (.A(net637),
    .B(net634),
    .C(net628),
    .Y(_0956_));
 sg13g2_a221oi_1 _2881_ (.B2(_0956_),
    .C1(net607),
    .B1(_0714_),
    .A1(net611),
    .Y(_0967_),
    .A2(_0659_));
 sg13g2_xnor2_1 _2882_ (.Y(_0978_),
    .A(net556),
    .B(_0967_));
 sg13g2_xnor2_1 _2883_ (.Y(_0989_),
    .A(net623),
    .B(_0967_));
 sg13g2_nand2_2 _2884_ (.Y(_0999_),
    .A(net652),
    .B(_0989_));
 sg13g2_xor2_1 _2885_ (.B(net643),
    .A(net647),
    .X(_1010_));
 sg13g2_xnor2_1 _2886_ (.Y(_1021_),
    .A(net649),
    .B(net643));
 sg13g2_mux2_1 _2887_ (.A0(_2668_),
    .A1(_1021_),
    .S(_0681_),
    .X(_1032_));
 sg13g2_mux2_1 _2888_ (.A0(net646),
    .A1(_1010_),
    .S(_0681_),
    .X(_1043_));
 sg13g2_a221oi_1 _2889_ (.B2(net547),
    .C1(net607),
    .B1(_0714_),
    .A1(net611),
    .Y(_1054_),
    .A2(_0659_));
 sg13g2_xor2_1 _2890_ (.B(_1054_),
    .A(net628),
    .X(_1065_));
 sg13g2_xnor2_1 _2891_ (.Y(_1076_),
    .A(net628),
    .B(_1054_));
 sg13g2_nor2_2 _2892_ (.A(_1032_),
    .B(net508),
    .Y(_1087_));
 sg13g2_nor2_2 _2893_ (.A(net567),
    .B(_0538_),
    .Y(_1098_));
 sg13g2_nand2_2 _2894_ (.Y(_1109_),
    .A(net563),
    .B(_0549_));
 sg13g2_nor2_1 _2895_ (.A(net567),
    .B(net589),
    .Y(_1120_));
 sg13g2_and2_1 _2896_ (.A(net582),
    .B(net587),
    .X(_1131_));
 sg13g2_nand2_2 _2897_ (.Y(_1141_),
    .A(net582),
    .B(net590));
 sg13g2_nand3_1 _2898_ (.B(net580),
    .C(net591),
    .A(net576),
    .Y(_1152_));
 sg13g2_and4_1 _2899_ (.A(net572),
    .B(net579),
    .C(net582),
    .D(net587),
    .X(_1163_));
 sg13g2_nand4_1 _2900_ (.B(net579),
    .C(net582),
    .A(net572),
    .Y(_1174_),
    .D(net587));
 sg13g2_nand2_2 _2901_ (.Y(_1185_),
    .A(net562),
    .B(_1174_));
 sg13g2_nor2_1 _2902_ (.A(net568),
    .B(_1163_),
    .Y(_1196_));
 sg13g2_nand2_1 _2903_ (.Y(_1207_),
    .A(_2613_),
    .B(_2624_));
 sg13g2_nor2_1 _2904_ (.A(net598),
    .B(net601),
    .Y(_1218_));
 sg13g2_nand2_2 _2905_ (.Y(_1229_),
    .A(_2624_),
    .B(_2635_));
 sg13g2_nor3_2 _2906_ (.A(net596),
    .B(net599),
    .C(net603),
    .Y(_1240_));
 sg13g2_or3_1 _2907_ (.A(net595),
    .B(net598),
    .C(net601),
    .X(_1251_));
 sg13g2_nor2_2 _2908_ (.A(net594),
    .B(net596),
    .Y(_1262_));
 sg13g2_nand2_2 _2909_ (.Y(_1273_),
    .A(net560),
    .B(_2613_));
 sg13g2_or4_1 _2910_ (.A(net593),
    .B(net596),
    .C(net599),
    .D(net603),
    .X(_1284_));
 sg13g2_a221oi_1 _2911_ (.B2(_1284_),
    .C1(net567),
    .B1(_1131_),
    .A1(net589),
    .Y(_1295_),
    .A2(_0538_));
 sg13g2_a21oi_2 _2912_ (.B1(net570),
    .Y(_1306_),
    .A2(\flag.flag_abrosexual_inst.pix_y[6] ),
    .A1(net576));
 sg13g2_nand2_2 _2913_ (.Y(_1317_),
    .A(net563),
    .B(_0505_));
 sg13g2_nor2_1 _2914_ (.A(_1141_),
    .B(net545),
    .Y(_1328_));
 sg13g2_or3_1 _2915_ (.A(net580),
    .B(_1295_),
    .C(_1328_),
    .X(_1339_));
 sg13g2_o21ai_1 _2916_ (.B1(net580),
    .Y(_1350_),
    .A1(_1295_),
    .A2(_1328_));
 sg13g2_and2_1 _2917_ (.A(_1339_),
    .B(_1350_),
    .X(_1361_));
 sg13g2_nand3_1 _2918_ (.B(_1339_),
    .C(_1350_),
    .A(net604),
    .Y(_1372_));
 sg13g2_nand3_1 _2919_ (.B(_1087_),
    .C(net462),
    .A(net604),
    .Y(_1383_));
 sg13g2_xor2_1 _2920_ (.B(_1372_),
    .A(_1087_),
    .X(_1394_));
 sg13g2_xor2_1 _2921_ (.B(_1394_),
    .A(_0999_),
    .X(_1405_));
 sg13g2_nor2_1 _2922_ (.A(net513),
    .B(_0868_),
    .Y(_1416_));
 sg13g2_nor2_2 _2923_ (.A(net558),
    .B(net557),
    .Y(_1427_));
 sg13g2_nor2_2 _2924_ (.A(net547),
    .B(_1427_),
    .Y(_1438_));
 sg13g2_a22oi_1 _2925_ (.Y(_1449_),
    .B1(_1416_),
    .B2(_1438_),
    .A2(_1405_),
    .A1(_0901_));
 sg13g2_nand2_2 _2926_ (.Y(_1460_),
    .A(net515),
    .B(net510));
 sg13g2_nor2_1 _2927_ (.A(net513),
    .B(_1460_),
    .Y(_1471_));
 sg13g2_and3_1 _2928_ (.X(_1482_),
    .A(net578),
    .B(net584),
    .C(net588));
 sg13g2_nand2_1 _2929_ (.Y(_1493_),
    .A(net579),
    .B(_1131_));
 sg13g2_a21o_1 _2930_ (.A2(_1482_),
    .A1(_1284_),
    .B1(net573),
    .X(_1504_));
 sg13g2_a21oi_1 _2931_ (.A1(net589),
    .A2(_1284_),
    .Y(_1515_),
    .B1(net567));
 sg13g2_o21ai_1 _2932_ (.B1(_1504_),
    .Y(_1526_),
    .A1(_1098_),
    .A2(_1515_));
 sg13g2_nor2_2 _2933_ (.A(net564),
    .B(net573),
    .Y(_1537_));
 sg13g2_nand2_1 _2934_ (.Y(_1548_),
    .A(net567),
    .B(_2569_));
 sg13g2_a21oi_2 _2935_ (.B1(_1163_),
    .Y(_1559_),
    .A2(_1537_),
    .A1(_1493_));
 sg13g2_and2_1 _2936_ (.A(_1526_),
    .B(_1559_),
    .X(_1570_));
 sg13g2_nand2_2 _2937_ (.Y(_1581_),
    .A(_1526_),
    .B(_1559_));
 sg13g2_nand3_1 _2938_ (.B(_1526_),
    .C(_1559_),
    .A(net604),
    .Y(_1592_));
 sg13g2_nand2_2 _2939_ (.Y(_1603_),
    .A(net515),
    .B(_1065_));
 sg13g2_nor2_1 _2940_ (.A(_0813_),
    .B(net508),
    .Y(_1614_));
 sg13g2_nor4_1 _2941_ (.A(net514),
    .B(_0813_),
    .C(_0868_),
    .D(net508),
    .Y(_1625_));
 sg13g2_nand4_1 _2942_ (.B(_0824_),
    .C(net511),
    .A(net515),
    .Y(_1636_),
    .D(_1065_));
 sg13g2_a22oi_1 _2943_ (.Y(_1647_),
    .B1(_1065_),
    .B2(_0824_),
    .A2(net511),
    .A1(net515));
 sg13g2_or3_1 _2944_ (.A(_1592_),
    .B(_1625_),
    .C(_1647_),
    .X(_1657_));
 sg13g2_o21ai_1 _2945_ (.B1(_1592_),
    .Y(_1668_),
    .A1(_1625_),
    .A2(_1647_));
 sg13g2_and3_1 _2946_ (.X(_1679_),
    .A(_1471_),
    .B(_1657_),
    .C(_1668_));
 sg13g2_nand3_1 _2947_ (.B(_1657_),
    .C(_1668_),
    .A(_1471_),
    .Y(_1690_));
 sg13g2_a21oi_1 _2948_ (.A1(_1657_),
    .A2(_1668_),
    .Y(_1701_),
    .B1(_1471_));
 sg13g2_a21o_1 _2949_ (.A2(_1668_),
    .A1(_1657_),
    .B1(_1471_),
    .X(_1712_));
 sg13g2_nor2_1 _2950_ (.A(net623),
    .B(net554),
    .Y(_1723_));
 sg13g2_nor2_2 _2951_ (.A(_2712_),
    .B(net617),
    .Y(_1734_));
 sg13g2_or2_1 _2952_ (.X(_1744_),
    .B(_1734_),
    .A(_1723_));
 sg13g2_nor2_2 _2953_ (.A(net614),
    .B(net607),
    .Y(_1755_));
 sg13g2_nand2_2 _2954_ (.Y(_1766_),
    .A(net552),
    .B(_2745_));
 sg13g2_a21oi_1 _2955_ (.A1(_0714_),
    .A2(_0956_),
    .Y(_1777_),
    .B1(_2712_));
 sg13g2_xnor2_1 _2956_ (.Y(_1788_),
    .A(net617),
    .B(_1777_));
 sg13g2_a22oi_1 _2957_ (.Y(_1799_),
    .B1(_1788_),
    .B2(_0681_),
    .A2(_1766_),
    .A1(_1744_));
 sg13g2_nand2_2 _2958_ (.Y(_1810_),
    .A(net652),
    .B(net461));
 sg13g2_nand2_2 _2959_ (.Y(_1821_),
    .A(_0989_),
    .B(net509));
 sg13g2_a21oi_2 _2960_ (.B1(net599),
    .Y(_1832_),
    .A2(_1174_),
    .A1(net562));
 sg13g2_nor3_1 _2961_ (.A(net566),
    .B(_2624_),
    .C(_1163_),
    .Y(_1843_));
 sg13g2_nor2_2 _2962_ (.A(_1832_),
    .B(_1843_),
    .Y(_1853_));
 sg13g2_o21ai_1 _2963_ (.B1(net600),
    .Y(_1864_),
    .A1(_1832_),
    .A2(_1843_));
 sg13g2_nand2_2 _2964_ (.Y(_1875_),
    .A(net603),
    .B(_1853_));
 sg13g2_and2_1 _2965_ (.A(net533),
    .B(net507),
    .X(_1886_));
 sg13g2_nand2_2 _2966_ (.Y(_1897_),
    .A(net533),
    .B(net507));
 sg13g2_nand4_1 _2967_ (.B(_1339_),
    .C(_1350_),
    .A(net533),
    .Y(_1908_),
    .D(net507));
 sg13g2_xor2_1 _2968_ (.B(_1908_),
    .A(_1821_),
    .X(_1917_));
 sg13g2_nand2b_1 _2969_ (.Y(_1922_),
    .B(_1917_),
    .A_N(_1810_));
 sg13g2_xnor2_1 _2970_ (.Y(_1927_),
    .A(_1810_),
    .B(_1917_));
 sg13g2_xor2_1 _2971_ (.B(_1917_),
    .A(_1810_),
    .X(_1934_));
 sg13g2_nor3_1 _2972_ (.A(_1679_),
    .B(_1701_),
    .C(_1934_),
    .Y(_1943_));
 sg13g2_a21oi_1 _2973_ (.A1(_1690_),
    .A2(_1712_),
    .Y(_1950_),
    .B1(_1927_));
 sg13g2_o21ai_1 _2974_ (.B1(_1927_),
    .Y(_1959_),
    .A1(_1679_),
    .A2(_1701_));
 sg13g2_nand3_1 _2975_ (.B(_1712_),
    .C(_1934_),
    .A(_1690_),
    .Y(_1970_));
 sg13g2_nor3_2 _2976_ (.A(_1449_),
    .B(_1943_),
    .C(_1950_),
    .Y(_1980_));
 sg13g2_or3_1 _2977_ (.A(_1449_),
    .B(_1943_),
    .C(_1950_),
    .X(_1990_));
 sg13g2_and3_1 _2978_ (.X(_2000_),
    .A(_1449_),
    .B(_1959_),
    .C(_1970_));
 sg13g2_o21ai_1 _2979_ (.B1(_1449_),
    .Y(_2009_),
    .A1(_1943_),
    .A2(_1950_));
 sg13g2_nor2_2 _2980_ (.A(net588),
    .B(net593),
    .Y(_2019_));
 sg13g2_nand2_1 _2981_ (.Y(_2023_),
    .A(_1240_),
    .B(_2019_));
 sg13g2_nand2_1 _2982_ (.Y(_2024_),
    .A(_1515_),
    .B(_2023_));
 sg13g2_nand2_1 _2983_ (.Y(_2025_),
    .A(net589),
    .B(_1109_));
 sg13g2_a22oi_1 _2984_ (.Y(_2026_),
    .B1(_1515_),
    .B2(_2023_),
    .A2(_1109_),
    .A1(net589));
 sg13g2_nand2_2 _2985_ (.Y(_2027_),
    .A(_2024_),
    .B(_2025_));
 sg13g2_nand3_1 _2986_ (.B(net507),
    .C(net505),
    .A(net533),
    .Y(_2028_));
 sg13g2_a21o_1 _2987_ (.A2(_1284_),
    .A1(net589),
    .B1(net584),
    .X(_2029_));
 sg13g2_or2_1 _2988_ (.X(_2030_),
    .B(net587),
    .A(net582));
 sg13g2_nand2_1 _2989_ (.Y(_2031_),
    .A(_1141_),
    .B(_2030_));
 sg13g2_and2_1 _2990_ (.A(_0494_),
    .B(net544),
    .X(_2032_));
 sg13g2_nor2_1 _2991_ (.A(net568),
    .B(_2032_),
    .Y(_2033_));
 sg13g2_a22oi_1 _2992_ (.Y(_2034_),
    .B1(_2031_),
    .B2(_1109_),
    .A2(_2029_),
    .A1(_1295_));
 sg13g2_o21ai_1 _2993_ (.B1(net596),
    .Y(_2035_),
    .A1(net566),
    .A2(_1163_));
 sg13g2_o21ai_1 _2994_ (.B1(net597),
    .Y(_2036_),
    .A1(net599),
    .A2(net601));
 sg13g2_nand2_1 _2995_ (.Y(_2037_),
    .A(_1251_),
    .B(_2036_));
 sg13g2_nor2_1 _2996_ (.A(net536),
    .B(_2037_),
    .Y(_2038_));
 sg13g2_a21oi_2 _2997_ (.B1(_2038_),
    .Y(_2039_),
    .A2(net536),
    .A1(net596));
 sg13g2_o21ai_1 _2998_ (.B1(_2035_),
    .Y(_2040_),
    .A1(net536),
    .A2(_2037_));
 sg13g2_nand2_2 _2999_ (.Y(_2041_),
    .A(net503),
    .B(_2040_));
 sg13g2_nand3_1 _3000_ (.B(_1864_),
    .C(net504),
    .A(_1229_),
    .Y(_2042_));
 sg13g2_inv_1 _3001_ (.Y(_2043_),
    .A(_2042_));
 sg13g2_nand2_2 _3002_ (.Y(_2044_),
    .A(net505),
    .B(net501));
 sg13g2_or2_1 _3003_ (.X(_2045_),
    .B(_2044_),
    .A(_2042_));
 sg13g2_o21ai_1 _3004_ (.B1(net592),
    .Y(_2046_),
    .A1(net566),
    .A2(_1163_));
 sg13g2_xnor2_1 _3005_ (.Y(_2047_),
    .A(net560),
    .B(_1240_));
 sg13g2_o21ai_1 _3006_ (.B1(_2046_),
    .Y(_2048_),
    .A1(net536),
    .A2(_2047_));
 sg13g2_inv_4 _3007_ (.A(net500),
    .Y(_2049_));
 sg13g2_and2_1 _3008_ (.A(_2042_),
    .B(_2044_),
    .X(_2050_));
 sg13g2_xor2_1 _3009_ (.B(_2044_),
    .A(_2042_),
    .X(_2051_));
 sg13g2_o21ai_1 _3010_ (.B1(_2045_),
    .Y(_2052_),
    .A1(_2049_),
    .A2(_2050_));
 sg13g2_o21ai_1 _3011_ (.B1(_1383_),
    .Y(_2053_),
    .A1(_0999_),
    .A2(_1394_));
 sg13g2_nor2b_1 _3012_ (.A(net460),
    .B_N(_2053_),
    .Y(_2054_));
 sg13g2_nand2b_1 _3013_ (.Y(_2055_),
    .B(net460),
    .A_N(_2053_));
 sg13g2_xor2_1 _3014_ (.B(_2053_),
    .A(net460),
    .X(_2056_));
 sg13g2_xnor2_1 _3015_ (.Y(_2057_),
    .A(_2052_),
    .B(_2056_));
 sg13g2_xor2_1 _3016_ (.B(_2056_),
    .A(_2052_),
    .X(_2058_));
 sg13g2_nor3_1 _3017_ (.A(_1980_),
    .B(_2000_),
    .C(_2058_),
    .Y(_2059_));
 sg13g2_a21oi_1 _3018_ (.A1(_2009_),
    .A2(_2057_),
    .Y(_2060_),
    .B1(_1980_));
 sg13g2_o21ai_1 _3019_ (.B1(_1690_),
    .Y(_2061_),
    .A1(_1701_),
    .A2(_1934_));
 sg13g2_o21ai_1 _3020_ (.B1(_1636_),
    .Y(_2062_),
    .A1(_1592_),
    .A2(_1647_));
 sg13g2_nand4_1 _3021_ (.B(_1526_),
    .C(_1559_),
    .A(_1229_),
    .Y(_2063_),
    .D(_1864_));
 sg13g2_nor2_1 _3022_ (.A(_0978_),
    .B(_1076_),
    .Y(_2064_));
 sg13g2_nand2_1 _3023_ (.Y(_2065_),
    .A(net511),
    .B(_1065_));
 sg13g2_nand2_1 _3024_ (.Y(_2066_),
    .A(net512),
    .B(_0989_));
 sg13g2_nor4_1 _3025_ (.A(_0813_),
    .B(_0868_),
    .C(_0978_),
    .D(_1076_),
    .Y(_2067_));
 sg13g2_a22oi_1 _3026_ (.Y(_2068_),
    .B1(_1065_),
    .B2(net511),
    .A2(_0989_),
    .A1(_0824_));
 sg13g2_or3_1 _3027_ (.A(_2063_),
    .B(_2067_),
    .C(_2068_),
    .X(_2069_));
 sg13g2_o21ai_1 _3028_ (.B1(_2063_),
    .Y(_2070_),
    .A1(_2067_),
    .A2(_2068_));
 sg13g2_and3_1 _3029_ (.X(_2071_),
    .A(_2062_),
    .B(_2069_),
    .C(_2070_));
 sg13g2_a21oi_1 _3030_ (.A1(_2069_),
    .A2(_2070_),
    .Y(_2072_),
    .B1(_2062_));
 sg13g2_nand2_2 _3031_ (.Y(_2073_),
    .A(net463),
    .B(net502));
 sg13g2_nand2_2 _3032_ (.Y(_2074_),
    .A(_1043_),
    .B(net461));
 sg13g2_or2_1 _3033_ (.X(_2075_),
    .B(_2074_),
    .A(_2073_));
 sg13g2_xnor2_1 _3034_ (.Y(_2076_),
    .A(_2073_),
    .B(_2074_));
 sg13g2_or3_1 _3035_ (.A(_2071_),
    .B(_2072_),
    .C(_2076_),
    .X(_2077_));
 sg13g2_o21ai_1 _3036_ (.B1(_2076_),
    .Y(_2078_),
    .A1(_2071_),
    .A2(_2072_));
 sg13g2_and3_1 _3037_ (.X(_2079_),
    .A(_2061_),
    .B(_2077_),
    .C(_2078_));
 sg13g2_nand3_1 _3038_ (.B(_2077_),
    .C(_2078_),
    .A(_2061_),
    .Y(_2080_));
 sg13g2_a21oi_1 _3039_ (.A1(_2077_),
    .A2(_2078_),
    .Y(_2081_),
    .B1(_2061_));
 sg13g2_a21o_1 _3040_ (.A2(_2078_),
    .A1(_2077_),
    .B1(_2061_),
    .X(_2082_));
 sg13g2_o21ai_1 _3041_ (.B1(_1922_),
    .Y(_2083_),
    .A1(_1821_),
    .A2(_1908_));
 sg13g2_nor2_1 _3042_ (.A(_2027_),
    .B(net499),
    .Y(_2084_));
 sg13g2_xor2_1 _3043_ (.B(_2084_),
    .A(_2083_),
    .X(_2085_));
 sg13g2_xnor2_1 _3044_ (.Y(_2086_),
    .A(_2083_),
    .B(_2084_));
 sg13g2_nor3_1 _3045_ (.A(_2079_),
    .B(_2081_),
    .C(_2086_),
    .Y(_2087_));
 sg13g2_nand3_1 _3046_ (.B(_2082_),
    .C(_2085_),
    .A(_2080_),
    .Y(_2088_));
 sg13g2_a21oi_1 _3047_ (.A1(_2080_),
    .A2(_2082_),
    .Y(_2089_),
    .B1(_2085_));
 sg13g2_o21ai_1 _3048_ (.B1(_2086_),
    .Y(_2090_),
    .A1(_2079_),
    .A2(_2081_));
 sg13g2_nor3_1 _3049_ (.A(_2060_),
    .B(_2087_),
    .C(_2089_),
    .Y(_2091_));
 sg13g2_nand3b_1 _3050_ (.B(_2088_),
    .C(_2090_),
    .Y(_2092_),
    .A_N(_2060_));
 sg13g2_a221oi_1 _3051_ (.B2(_2090_),
    .C1(_1980_),
    .B1(_2088_),
    .A1(_2009_),
    .Y(_2093_),
    .A2(_2057_));
 sg13g2_o21ai_1 _3052_ (.B1(_2060_),
    .Y(_2094_),
    .A1(_2087_),
    .A2(_2089_));
 sg13g2_o21ai_1 _3053_ (.B1(_2045_),
    .Y(_2095_),
    .A1(_1372_),
    .A2(_2050_));
 sg13g2_and3_2 _3054_ (.X(_2096_),
    .A(net533),
    .B(net507),
    .C(net501));
 sg13g2_nand3_1 _3055_ (.B(net507),
    .C(net501),
    .A(net533),
    .Y(_2097_));
 sg13g2_nand2_2 _3056_ (.Y(_2098_),
    .A(net462),
    .B(net503));
 sg13g2_or2_1 _3057_ (.X(_2099_),
    .B(net460),
    .A(_1908_));
 sg13g2_and2_1 _3058_ (.A(_1908_),
    .B(_2041_),
    .X(_2100_));
 sg13g2_xor2_1 _3059_ (.B(_2041_),
    .A(_1908_),
    .X(_2101_));
 sg13g2_xnor2_1 _3060_ (.Y(_2102_),
    .A(_1592_),
    .B(_2101_));
 sg13g2_nand2_1 _3061_ (.Y(_2103_),
    .A(_2095_),
    .B(_2102_));
 sg13g2_xnor2_1 _3062_ (.Y(_2104_),
    .A(_2095_),
    .B(_2102_));
 sg13g2_nand2_1 _3063_ (.Y(_2105_),
    .A(_0989_),
    .B(net461));
 sg13g2_xor2_1 _3064_ (.B(_1821_),
    .A(_1810_),
    .X(_2106_));
 sg13g2_nand2_1 _3065_ (.Y(_2107_),
    .A(_1614_),
    .B(_2106_));
 sg13g2_xnor2_1 _3066_ (.Y(_2108_),
    .A(_1614_),
    .B(_2106_));
 sg13g2_o21ai_1 _3067_ (.B1(_2103_),
    .Y(_2109_),
    .A1(_2104_),
    .A2(_2108_));
 sg13g2_a21oi_2 _3068_ (.B1(_2054_),
    .Y(_2110_),
    .A2(_2055_),
    .A1(_2052_));
 sg13g2_o21ai_1 _3069_ (.B1(_2099_),
    .Y(_2111_),
    .A1(_1592_),
    .A2(_2100_));
 sg13g2_and2_1 _3070_ (.A(net463),
    .B(_1570_),
    .X(_2112_));
 sg13g2_xor2_1 _3071_ (.B(_2073_),
    .A(_2063_),
    .X(_2113_));
 sg13g2_nand2_1 _3072_ (.Y(_2114_),
    .A(_2111_),
    .B(_2113_));
 sg13g2_xnor2_1 _3073_ (.Y(_2115_),
    .A(_2111_),
    .B(_2113_));
 sg13g2_a221oi_1 _3074_ (.B2(_0681_),
    .C1(net513),
    .B1(_1788_),
    .A1(_1744_),
    .Y(_2116_),
    .A2(_1766_));
 sg13g2_xor2_1 _3075_ (.B(_2074_),
    .A(_2066_),
    .X(_2117_));
 sg13g2_nand2b_1 _3076_ (.Y(_2118_),
    .B(_2117_),
    .A_N(_2065_));
 sg13g2_xor2_1 _3077_ (.B(_2117_),
    .A(_2065_),
    .X(_2119_));
 sg13g2_xor2_1 _3078_ (.B(_2119_),
    .A(_2115_),
    .X(_2120_));
 sg13g2_nor2b_1 _3079_ (.A(_2110_),
    .B_N(_2120_),
    .Y(_2121_));
 sg13g2_xnor2_1 _3080_ (.Y(_2122_),
    .A(_2110_),
    .B(_2120_));
 sg13g2_xor2_1 _3081_ (.B(_2122_),
    .A(_2109_),
    .X(_2123_));
 sg13g2_xnor2_1 _3082_ (.Y(_2124_),
    .A(_2109_),
    .B(_2122_));
 sg13g2_nor3_1 _3083_ (.A(_2091_),
    .B(_2093_),
    .C(_2124_),
    .Y(_2125_));
 sg13g2_nor2_1 _3084_ (.A(_2091_),
    .B(_2125_),
    .Y(_2126_));
 sg13g2_nand2_1 _3085_ (.Y(_2127_),
    .A(_2080_),
    .B(_2088_));
 sg13g2_nand2b_1 _3086_ (.Y(_2128_),
    .B(_2077_),
    .A_N(_2071_));
 sg13g2_nand2_1 _3087_ (.Y(_2129_),
    .A(net463),
    .B(net499));
 sg13g2_inv_1 _3088_ (.Y(_2130_),
    .A(_2129_));
 sg13g2_nor2b_1 _3089_ (.A(_2067_),
    .B_N(_2069_),
    .Y(_2131_));
 sg13g2_nand2_1 _3090_ (.Y(_2132_),
    .A(_1570_),
    .B(net502));
 sg13g2_nor2_1 _3091_ (.A(_0868_),
    .B(_0978_),
    .Y(_2133_));
 sg13g2_nand2_1 _3092_ (.Y(_2134_),
    .A(_2116_),
    .B(_2133_));
 sg13g2_xnor2_1 _3093_ (.Y(_2135_),
    .A(_2116_),
    .B(_2133_));
 sg13g2_xnor2_1 _3094_ (.Y(_2136_),
    .A(_2132_),
    .B(_2135_));
 sg13g2_nor2_1 _3095_ (.A(_2131_),
    .B(_2136_),
    .Y(_2137_));
 sg13g2_xor2_1 _3096_ (.B(_2136_),
    .A(_2131_),
    .X(_2138_));
 sg13g2_xnor2_1 _3097_ (.Y(_2139_),
    .A(_2129_),
    .B(_2138_));
 sg13g2_nand2_1 _3098_ (.Y(_2140_),
    .A(_2128_),
    .B(_2139_));
 sg13g2_xnor2_1 _3099_ (.Y(_2141_),
    .A(_2128_),
    .B(_2139_));
 sg13g2_nand2_2 _3100_ (.Y(_2142_),
    .A(net503),
    .B(net500));
 sg13g2_mux2_1 _3101_ (.A0(net499),
    .A1(_2129_),
    .S(_2075_),
    .X(_2143_));
 sg13g2_or2_1 _3102_ (.X(_2144_),
    .B(_2143_),
    .A(_2142_));
 sg13g2_xnor2_1 _3103_ (.Y(_2145_),
    .A(_2142_),
    .B(_2143_));
 sg13g2_xor2_1 _3104_ (.B(_2145_),
    .A(_2141_),
    .X(_2146_));
 sg13g2_nand2_1 _3105_ (.Y(_2147_),
    .A(_2127_),
    .B(_2146_));
 sg13g2_xnor2_1 _3106_ (.Y(_2148_),
    .A(_2127_),
    .B(_2146_));
 sg13g2_o21ai_1 _3107_ (.B1(_2114_),
    .Y(_2149_),
    .A1(_2115_),
    .A2(_2119_));
 sg13g2_nand3_1 _3108_ (.B(_1908_),
    .C(net502),
    .A(_1570_),
    .Y(_2150_));
 sg13g2_xnor2_1 _3109_ (.Y(_2151_),
    .A(_1603_),
    .B(_2135_));
 sg13g2_nor2_1 _3110_ (.A(_2150_),
    .B(_2151_),
    .Y(_2152_));
 sg13g2_xnor2_1 _3111_ (.Y(_2153_),
    .A(_2150_),
    .B(_2151_));
 sg13g2_and2_1 _3112_ (.A(net505),
    .B(net500),
    .X(_2154_));
 sg13g2_nand2_1 _3113_ (.Y(_2155_),
    .A(net505),
    .B(net500));
 sg13g2_o21ai_1 _3114_ (.B1(net505),
    .Y(_2156_),
    .A1(net499),
    .A2(_2083_));
 sg13g2_nor2_1 _3115_ (.A(_2153_),
    .B(_2156_),
    .Y(_2157_));
 sg13g2_xor2_1 _3116_ (.B(_2156_),
    .A(_2153_),
    .X(_2158_));
 sg13g2_xnor2_1 _3117_ (.Y(_2159_),
    .A(_2149_),
    .B(_2158_));
 sg13g2_xor2_1 _3118_ (.B(_2159_),
    .A(_2148_),
    .X(_2160_));
 sg13g2_nand2b_1 _3119_ (.Y(_2161_),
    .B(_2160_),
    .A_N(_2126_));
 sg13g2_xor2_1 _3120_ (.B(_2160_),
    .A(_2126_),
    .X(_2162_));
 sg13g2_a21oi_1 _3121_ (.A1(_2109_),
    .A2(_2122_),
    .Y(_2163_),
    .B1(_2121_));
 sg13g2_o21ai_1 _3122_ (.B1(_2118_),
    .Y(_2164_),
    .A1(_2066_),
    .A2(_2074_));
 sg13g2_nand2b_1 _3123_ (.Y(_2165_),
    .B(_2164_),
    .A_N(_2163_));
 sg13g2_xor2_1 _3124_ (.B(_2164_),
    .A(_2163_),
    .X(_2166_));
 sg13g2_xnor2_1 _3125_ (.Y(_2167_),
    .A(_1603_),
    .B(_2166_));
 sg13g2_o21ai_1 _3126_ (.B1(_2161_),
    .Y(_2168_),
    .A1(_2162_),
    .A2(_2167_));
 sg13g2_o21ai_1 _3127_ (.B1(_2147_),
    .Y(_2169_),
    .A1(_2148_),
    .A2(_2159_));
 sg13g2_o21ai_1 _3128_ (.B1(_2140_),
    .Y(_2170_),
    .A1(_2141_),
    .A2(_2145_));
 sg13g2_nand2_2 _3129_ (.Y(_2171_),
    .A(net506),
    .B(net504));
 sg13g2_nand2_2 _3130_ (.Y(_2172_),
    .A(_1570_),
    .B(net499));
 sg13g2_nand2_2 _3131_ (.Y(_2173_),
    .A(net462),
    .B(net506));
 sg13g2_xor2_1 _3132_ (.B(_2173_),
    .A(net503),
    .X(_2174_));
 sg13g2_or2_1 _3133_ (.X(_2175_),
    .B(_2174_),
    .A(_2172_));
 sg13g2_xor2_1 _3134_ (.B(_2174_),
    .A(_2172_),
    .X(_2176_));
 sg13g2_nand2b_1 _3135_ (.Y(_2177_),
    .B(_2176_),
    .A_N(_2171_));
 sg13g2_xnor2_1 _3136_ (.Y(_2178_),
    .A(_2171_),
    .B(_2176_));
 sg13g2_a21oi_1 _3137_ (.A1(_2130_),
    .A2(_2138_),
    .Y(_2179_),
    .B1(_2137_));
 sg13g2_o21ai_1 _3138_ (.B1(_2134_),
    .Y(_2180_),
    .A1(_2132_),
    .A2(_2135_));
 sg13g2_nand2_2 _3139_ (.Y(_2181_),
    .A(net511),
    .B(net461));
 sg13g2_or2_1 _3140_ (.X(_2182_),
    .B(_2181_),
    .A(_2172_));
 sg13g2_xor2_1 _3141_ (.B(_2181_),
    .A(_2172_),
    .X(_2183_));
 sg13g2_nand2_1 _3142_ (.Y(_2184_),
    .A(_2180_),
    .B(_2183_));
 sg13g2_xnor2_1 _3143_ (.Y(_2185_),
    .A(_2180_),
    .B(_2183_));
 sg13g2_xor2_1 _3144_ (.B(_2185_),
    .A(_2173_),
    .X(_2186_));
 sg13g2_nor2b_1 _3145_ (.A(_2179_),
    .B_N(_2186_),
    .Y(_2187_));
 sg13g2_xnor2_1 _3146_ (.Y(_2188_),
    .A(_2179_),
    .B(_2186_));
 sg13g2_xnor2_1 _3147_ (.Y(_2189_),
    .A(_2178_),
    .B(_2188_));
 sg13g2_nand2b_1 _3148_ (.Y(_2190_),
    .B(_2170_),
    .A_N(_2189_));
 sg13g2_xor2_1 _3149_ (.B(_2189_),
    .A(_2170_),
    .X(_2191_));
 sg13g2_a21oi_1 _3150_ (.A1(_2096_),
    .A2(_2112_),
    .Y(_2192_),
    .B1(_2152_));
 sg13g2_o21ai_1 _3151_ (.B1(_2144_),
    .Y(_2193_),
    .A1(_2049_),
    .A2(_2075_));
 sg13g2_nand2_2 _3152_ (.Y(_2194_),
    .A(net515),
    .B(_0989_));
 sg13g2_nand2_2 _3153_ (.Y(_2195_),
    .A(net515),
    .B(net461));
 sg13g2_nor2_1 _3154_ (.A(_1460_),
    .B(_2105_),
    .Y(_2196_));
 sg13g2_a21oi_1 _3155_ (.A1(_2181_),
    .A2(_2194_),
    .Y(_2197_),
    .B1(_2196_));
 sg13g2_xnor2_1 _3156_ (.Y(_2198_),
    .A(_1076_),
    .B(_2197_));
 sg13g2_nand2_1 _3157_ (.Y(_2199_),
    .A(_2193_),
    .B(_2198_));
 sg13g2_xnor2_1 _3158_ (.Y(_2200_),
    .A(_2193_),
    .B(_2198_));
 sg13g2_xnor2_1 _3159_ (.Y(_2201_),
    .A(_2192_),
    .B(_2200_));
 sg13g2_xor2_1 _3160_ (.B(_2201_),
    .A(_2191_),
    .X(_2202_));
 sg13g2_nand2_1 _3161_ (.Y(_2203_),
    .A(_2169_),
    .B(_2202_));
 sg13g2_xnor2_1 _3162_ (.Y(_2204_),
    .A(_2169_),
    .B(_2202_));
 sg13g2_a21oi_1 _3163_ (.A1(_2149_),
    .A2(_2158_),
    .Y(_2205_),
    .B1(_2157_));
 sg13g2_o21ai_1 _3164_ (.B1(_2134_),
    .Y(_2206_),
    .A1(_1603_),
    .A2(_2135_));
 sg13g2_nand2b_1 _3165_ (.Y(_2207_),
    .B(_2206_),
    .A_N(_2205_));
 sg13g2_xor2_1 _3166_ (.B(_2206_),
    .A(_2205_),
    .X(_2208_));
 sg13g2_xnor2_1 _3167_ (.Y(_2209_),
    .A(_2194_),
    .B(_2208_));
 sg13g2_xor2_1 _3168_ (.B(_2209_),
    .A(_2204_),
    .X(_2210_));
 sg13g2_nand2_1 _3169_ (.Y(_2211_),
    .A(_2168_),
    .B(_2210_));
 sg13g2_o21ai_1 _3170_ (.B1(_2165_),
    .Y(_2212_),
    .A1(_1603_),
    .A2(_2166_));
 sg13g2_xnor2_1 _3171_ (.Y(_2213_),
    .A(_2168_),
    .B(_2210_));
 sg13g2_nand2b_1 _3172_ (.Y(_2214_),
    .B(_2212_),
    .A_N(_2213_));
 sg13g2_o21ai_1 _3173_ (.B1(_2207_),
    .Y(_2215_),
    .A1(_2194_),
    .A2(_2208_));
 sg13g2_o21ai_1 _3174_ (.B1(_2203_),
    .Y(_2216_),
    .A1(_2204_),
    .A2(_2209_));
 sg13g2_o21ai_1 _3175_ (.B1(_2199_),
    .Y(_2217_),
    .A1(_2192_),
    .A2(_2200_));
 sg13g2_a21o_1 _3176_ (.A2(_2197_),
    .A1(_1065_),
    .B1(_2196_),
    .X(_2218_));
 sg13g2_xor2_1 _3177_ (.B(_2218_),
    .A(_2217_),
    .X(_2219_));
 sg13g2_nor2b_1 _3178_ (.A(_2195_),
    .B_N(_2219_),
    .Y(_2220_));
 sg13g2_xnor2_1 _3179_ (.Y(_2221_),
    .A(_2195_),
    .B(_2219_));
 sg13g2_o21ai_1 _3180_ (.B1(_2190_),
    .Y(_2222_),
    .A1(_2191_),
    .A2(_2201_));
 sg13g2_nor2_1 _3181_ (.A(_2177_),
    .B(_2195_),
    .Y(_2223_));
 sg13g2_xor2_1 _3182_ (.B(_2195_),
    .A(_2177_),
    .X(_2224_));
 sg13g2_a21oi_1 _3183_ (.A1(_2178_),
    .A2(_2188_),
    .Y(_2225_),
    .B1(_2187_));
 sg13g2_o21ai_1 _3184_ (.B1(_2175_),
    .Y(_2226_),
    .A1(_2027_),
    .A2(_2098_));
 sg13g2_nand2_1 _3185_ (.Y(_2227_),
    .A(_1570_),
    .B(net506));
 sg13g2_nand2_2 _3186_ (.Y(_2228_),
    .A(_1570_),
    .B(net503));
 sg13g2_xor2_1 _3187_ (.B(_2227_),
    .A(_2098_),
    .X(_2229_));
 sg13g2_nand2_1 _3188_ (.Y(_2230_),
    .A(_2226_),
    .B(_2229_));
 sg13g2_xnor2_1 _3189_ (.Y(_2231_),
    .A(_2226_),
    .B(_2229_));
 sg13g2_o21ai_1 _3190_ (.B1(_2184_),
    .Y(_2232_),
    .A1(_2173_),
    .A2(_2185_));
 sg13g2_or2_1 _3191_ (.X(_2233_),
    .B(_2182_),
    .A(_2027_));
 sg13g2_mux2_1 _3192_ (.A0(net506),
    .A1(_2227_),
    .S(_2182_),
    .X(_2234_));
 sg13g2_xor2_1 _3193_ (.B(_2234_),
    .A(_2098_),
    .X(_2235_));
 sg13g2_nand2_1 _3194_ (.Y(_2236_),
    .A(_2232_),
    .B(_2235_));
 sg13g2_xnor2_1 _3195_ (.Y(_2237_),
    .A(_2232_),
    .B(_2235_));
 sg13g2_xor2_1 _3196_ (.B(_2237_),
    .A(_2231_),
    .X(_2238_));
 sg13g2_nor2b_1 _3197_ (.A(_2225_),
    .B_N(_2238_),
    .Y(_2239_));
 sg13g2_xnor2_1 _3198_ (.Y(_2240_),
    .A(_2225_),
    .B(_2238_));
 sg13g2_xnor2_1 _3199_ (.Y(_2241_),
    .A(_2224_),
    .B(_2240_));
 sg13g2_nor2b_1 _3200_ (.A(_2241_),
    .B_N(_2222_),
    .Y(_2242_));
 sg13g2_xnor2_1 _3201_ (.Y(_2243_),
    .A(_2222_),
    .B(_2241_));
 sg13g2_xnor2_1 _3202_ (.Y(_2244_),
    .A(_2221_),
    .B(_2243_));
 sg13g2_nor2b_1 _3203_ (.A(_2244_),
    .B_N(_2216_),
    .Y(_2245_));
 sg13g2_xor2_1 _3204_ (.B(_2244_),
    .A(_2216_),
    .X(_2246_));
 sg13g2_inv_1 _3205_ (.Y(_2247_),
    .A(_2246_));
 sg13g2_xor2_1 _3206_ (.B(_2246_),
    .A(_2215_),
    .X(_2248_));
 sg13g2_and3_1 _3207_ (.X(_2249_),
    .A(_2211_),
    .B(_2214_),
    .C(_2248_));
 sg13g2_nand3_1 _3208_ (.B(_2214_),
    .C(_2248_),
    .A(_2211_),
    .Y(_2250_));
 sg13g2_xor2_1 _3209_ (.B(_2213_),
    .A(_2212_),
    .X(_2251_));
 sg13g2_nand2_2 _3210_ (.Y(_2252_),
    .A(net510),
    .B(net509));
 sg13g2_nor2_1 _3211_ (.A(net513),
    .B(_2252_),
    .Y(_2253_));
 sg13g2_nor2_1 _3212_ (.A(net559),
    .B(net514),
    .Y(_2254_));
 sg13g2_inv_1 _3213_ (.Y(_2255_),
    .A(_2254_));
 sg13g2_nor2_2 _3214_ (.A(net514),
    .B(_1032_),
    .Y(_2256_));
 sg13g2_nor2_2 _3215_ (.A(net559),
    .B(net508),
    .Y(_2257_));
 sg13g2_nand2_1 _3216_ (.Y(_2258_),
    .A(_1087_),
    .B(_2254_));
 sg13g2_xnor2_1 _3217_ (.Y(_2259_),
    .A(_2256_),
    .B(_2257_));
 sg13g2_nor3_1 _3218_ (.A(net513),
    .B(_2252_),
    .C(_2259_),
    .Y(_2260_));
 sg13g2_xnor2_1 _3219_ (.Y(_2261_),
    .A(_0890_),
    .B(_1405_));
 sg13g2_and2_1 _3220_ (.A(_2260_),
    .B(_2261_),
    .X(_2262_));
 sg13g2_or2_1 _3221_ (.X(_2263_),
    .B(_2261_),
    .A(_2260_));
 sg13g2_xnor2_1 _3222_ (.Y(_2264_),
    .A(_2260_),
    .B(_2261_));
 sg13g2_nand2_1 _3223_ (.Y(_2265_),
    .A(net501),
    .B(net500));
 sg13g2_nand3_1 _3224_ (.B(net507),
    .C(net500),
    .A(net533),
    .Y(_2266_));
 sg13g2_nand2b_1 _3225_ (.Y(_2267_),
    .B(net502),
    .A_N(_2266_));
 sg13g2_nor2_1 _3226_ (.A(_2097_),
    .B(_2155_),
    .Y(_2268_));
 sg13g2_and2_1 _3227_ (.A(net600),
    .B(net504),
    .X(_2269_));
 sg13g2_nand2_2 _3228_ (.Y(_2270_),
    .A(net603),
    .B(net504));
 sg13g2_a22oi_1 _3229_ (.Y(_2271_),
    .B1(_2265_),
    .B2(_2028_),
    .A2(_2154_),
    .A1(_2096_));
 sg13g2_a21oi_2 _3230_ (.B1(_2268_),
    .Y(_2272_),
    .A2(_2271_),
    .A1(_2269_));
 sg13g2_inv_1 _3231_ (.Y(_2273_),
    .A(_2272_));
 sg13g2_xnor2_1 _3232_ (.Y(_2274_),
    .A(net499),
    .B(_2051_));
 sg13g2_nor2_1 _3233_ (.A(_2258_),
    .B(_2274_),
    .Y(_2275_));
 sg13g2_xor2_1 _3234_ (.B(_2274_),
    .A(_2258_),
    .X(_2276_));
 sg13g2_xnor2_1 _3235_ (.Y(_2277_),
    .A(_2272_),
    .B(_2276_));
 sg13g2_a21oi_1 _3236_ (.A1(_2263_),
    .A2(_2277_),
    .Y(_2278_),
    .B1(_2262_));
 sg13g2_a21oi_1 _3237_ (.A1(_1990_),
    .A2(_2009_),
    .Y(_2279_),
    .B1(_2057_));
 sg13g2_o21ai_1 _3238_ (.B1(_2057_),
    .Y(_2280_),
    .A1(_1980_),
    .A2(_2000_));
 sg13g2_nand3_1 _3239_ (.B(_2009_),
    .C(_2058_),
    .A(_1990_),
    .Y(_2281_));
 sg13g2_nor3_1 _3240_ (.A(_2059_),
    .B(_2278_),
    .C(_2279_),
    .Y(_2282_));
 sg13g2_and3_1 _3241_ (.X(_2283_),
    .A(_2278_),
    .B(_2280_),
    .C(_2281_));
 sg13g2_o21ai_1 _3242_ (.B1(_2278_),
    .Y(_2284_),
    .A1(_2059_),
    .A2(_2279_));
 sg13g2_xnor2_1 _3243_ (.Y(_2285_),
    .A(_1372_),
    .B(_2051_));
 sg13g2_nor2b_1 _3244_ (.A(_2272_),
    .B_N(_2285_),
    .Y(_2286_));
 sg13g2_nand2b_1 _3245_ (.Y(_2287_),
    .B(_2257_),
    .A_N(_1821_));
 sg13g2_xnor2_1 _3246_ (.Y(_2288_),
    .A(_0999_),
    .B(_1087_));
 sg13g2_xnor2_1 _3247_ (.Y(_2289_),
    .A(_2272_),
    .B(_2285_));
 sg13g2_a21o_2 _3248_ (.A2(_2289_),
    .A1(_2288_),
    .B1(_2286_),
    .X(_2290_));
 sg13g2_a21oi_1 _3249_ (.A1(_2273_),
    .A2(_2276_),
    .Y(_2291_),
    .B1(_2275_));
 sg13g2_xor2_1 _3250_ (.B(_2108_),
    .A(_2104_),
    .X(_2292_));
 sg13g2_nor2b_1 _3251_ (.A(_2291_),
    .B_N(_2292_),
    .Y(_2293_));
 sg13g2_xnor2_1 _3252_ (.Y(_2294_),
    .A(_2291_),
    .B(_2292_));
 sg13g2_xor2_1 _3253_ (.B(_2294_),
    .A(_2290_),
    .X(_2295_));
 sg13g2_xnor2_1 _3254_ (.Y(_2296_),
    .A(_2290_),
    .B(_2294_));
 sg13g2_nand3b_1 _3255_ (.B(_2284_),
    .C(_2295_),
    .Y(_2297_),
    .A_N(_2282_));
 sg13g2_a21oi_2 _3256_ (.B1(_2282_),
    .Y(_2298_),
    .A2(_2295_),
    .A1(_2284_));
 sg13g2_a21oi_1 _3257_ (.A1(_2092_),
    .A2(_2094_),
    .Y(_2299_),
    .B1(_2123_));
 sg13g2_o21ai_1 _3258_ (.B1(_2123_),
    .Y(_2300_),
    .A1(_2091_),
    .A2(_2093_));
 sg13g2_nand3_1 _3259_ (.B(_2094_),
    .C(_2124_),
    .A(_2092_),
    .Y(_2301_));
 sg13g2_nor3_1 _3260_ (.A(_2125_),
    .B(_2298_),
    .C(_2299_),
    .Y(_2302_));
 sg13g2_or3_1 _3261_ (.A(_2125_),
    .B(_2298_),
    .C(_2299_),
    .X(_2303_));
 sg13g2_and3_1 _3262_ (.X(_2304_),
    .A(_2298_),
    .B(_2300_),
    .C(_2301_));
 sg13g2_o21ai_1 _3263_ (.B1(_2298_),
    .Y(_2305_),
    .A1(_2125_),
    .A2(_2299_));
 sg13g2_a21oi_1 _3264_ (.A1(_2290_),
    .A2(_2294_),
    .Y(_2306_),
    .B1(_2293_));
 sg13g2_o21ai_1 _3265_ (.B1(_2107_),
    .Y(_2307_),
    .A1(_1810_),
    .A2(_1821_));
 sg13g2_nand2b_1 _3266_ (.Y(_2308_),
    .B(_2307_),
    .A_N(_2306_));
 sg13g2_xor2_1 _3267_ (.B(_2307_),
    .A(_2306_),
    .X(_2309_));
 sg13g2_xnor2_1 _3268_ (.Y(_2310_),
    .A(_0780_),
    .B(_2309_));
 sg13g2_xnor2_1 _3269_ (.Y(_2311_),
    .A(_0791_),
    .B(_2309_));
 sg13g2_nor3_1 _3270_ (.A(_2302_),
    .B(_2304_),
    .C(_2311_),
    .Y(_2312_));
 sg13g2_nor2_1 _3271_ (.A(_2302_),
    .B(_2312_),
    .Y(_2313_));
 sg13g2_xnor2_1 _3272_ (.Y(_2314_),
    .A(_2162_),
    .B(_2167_));
 sg13g2_nor2_1 _3273_ (.A(_2313_),
    .B(_2314_),
    .Y(_2315_));
 sg13g2_o21ai_1 _3274_ (.B1(_2308_),
    .Y(_2316_),
    .A1(_0791_),
    .A2(_2309_));
 sg13g2_xor2_1 _3275_ (.B(_2314_),
    .A(_2313_),
    .X(_2317_));
 sg13g2_a21oi_1 _3276_ (.A1(_2316_),
    .A2(_2317_),
    .Y(_2318_),
    .B1(_2315_));
 sg13g2_nor2_1 _3277_ (.A(_2251_),
    .B(_2318_),
    .Y(_2319_));
 sg13g2_inv_1 _3278_ (.Y(_2320_),
    .A(_2319_));
 sg13g2_a21oi_1 _3279_ (.A1(_2211_),
    .A2(_2214_),
    .Y(_2321_),
    .B1(_2248_));
 sg13g2_o21ai_1 _3280_ (.B1(_2250_),
    .Y(_2322_),
    .A1(_2319_),
    .A2(_2321_));
 sg13g2_nor4_2 _3281_ (.A(net559),
    .B(net514),
    .C(_0868_),
    .Y(_2323_),
    .D(_1032_));
 sg13g2_a221oi_1 _3282_ (.B2(_2252_),
    .C1(_2323_),
    .B1(_0846_),
    .A1(_2646_),
    .Y(_2324_),
    .A2(net512));
 sg13g2_xor2_1 _3283_ (.B(_2259_),
    .A(_2253_),
    .X(_2325_));
 sg13g2_inv_1 _3284_ (.Y(_2326_),
    .A(_2325_));
 sg13g2_nand2_1 _3285_ (.Y(_2327_),
    .A(_2324_),
    .B(_2326_));
 sg13g2_xor2_1 _3286_ (.B(_2325_),
    .A(_2324_),
    .X(_2328_));
 sg13g2_xnor2_1 _3287_ (.Y(_2329_),
    .A(net560),
    .B(net537));
 sg13g2_xnor2_1 _3288_ (.Y(_2330_),
    .A(net592),
    .B(net536));
 sg13g2_nand2_2 _3289_ (.Y(_2331_),
    .A(net603),
    .B(net497));
 sg13g2_or2_1 _3290_ (.X(_2332_),
    .B(_2331_),
    .A(_2028_));
 sg13g2_xnor2_1 _3291_ (.Y(_2333_),
    .A(_2270_),
    .B(_2271_));
 sg13g2_nand2_1 _3292_ (.Y(_2334_),
    .A(_2323_),
    .B(_2333_));
 sg13g2_xnor2_1 _3293_ (.Y(_2335_),
    .A(_2323_),
    .B(_2333_));
 sg13g2_xnor2_1 _3294_ (.Y(_2336_),
    .A(_2332_),
    .B(_2335_));
 sg13g2_o21ai_1 _3295_ (.B1(_2327_),
    .Y(_2337_),
    .A1(_2328_),
    .A2(_2336_));
 sg13g2_xnor2_1 _3296_ (.Y(_2338_),
    .A(_2264_),
    .B(_2277_));
 sg13g2_nand2_1 _3297_ (.Y(_2339_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_xnor2_1 _3298_ (.Y(_2340_),
    .A(_2337_),
    .B(_2338_));
 sg13g2_nand2_2 _3299_ (.Y(_2341_),
    .A(net603),
    .B(net505));
 sg13g2_xnor2_1 _3300_ (.Y(_2342_),
    .A(_2039_),
    .B(_2266_));
 sg13g2_o21ai_1 _3301_ (.B1(_2267_),
    .Y(_2343_),
    .A1(_2341_),
    .A2(_2342_));
 sg13g2_and2_1 _3302_ (.A(_2333_),
    .B(_2343_),
    .X(_2344_));
 sg13g2_xor2_1 _3303_ (.B(_2343_),
    .A(_2333_),
    .X(_2345_));
 sg13g2_a21oi_1 _3304_ (.A1(_2257_),
    .A2(_2345_),
    .Y(_2346_),
    .B1(_2344_));
 sg13g2_o21ai_1 _3305_ (.B1(_2334_),
    .Y(_2347_),
    .A1(_2332_),
    .A2(_2335_));
 sg13g2_xnor2_1 _3306_ (.Y(_2348_),
    .A(_2288_),
    .B(_2289_));
 sg13g2_nand2b_1 _3307_ (.Y(_2349_),
    .B(_2347_),
    .A_N(_2348_));
 sg13g2_xor2_1 _3308_ (.B(_2348_),
    .A(_2347_),
    .X(_2350_));
 sg13g2_xnor2_1 _3309_ (.Y(_2351_),
    .A(_2346_),
    .B(_2350_));
 sg13g2_o21ai_1 _3310_ (.B1(_2339_),
    .Y(_2352_),
    .A1(_2340_),
    .A2(_2351_));
 sg13g2_o21ai_1 _3311_ (.B1(_2296_),
    .Y(_2353_),
    .A1(_2282_),
    .A2(_2283_));
 sg13g2_and3_1 _3312_ (.X(_2354_),
    .A(_2297_),
    .B(_2352_),
    .C(_2353_));
 sg13g2_nand3_1 _3313_ (.B(_2352_),
    .C(_2353_),
    .A(_2297_),
    .Y(_2355_));
 sg13g2_a21o_1 _3314_ (.A2(_2353_),
    .A1(_2297_),
    .B1(_2352_),
    .X(_2356_));
 sg13g2_o21ai_1 _3315_ (.B1(_2349_),
    .Y(_2357_),
    .A1(_2346_),
    .A2(_2350_));
 sg13g2_nand2b_1 _3316_ (.Y(_2358_),
    .B(_2357_),
    .A_N(_2287_));
 sg13g2_xor2_1 _3317_ (.B(_2357_),
    .A(_2287_),
    .X(_2359_));
 sg13g2_xor2_1 _3318_ (.B(_2359_),
    .A(_1460_),
    .X(_2360_));
 sg13g2_and3_2 _3319_ (.X(_2361_),
    .A(_2355_),
    .B(_2356_),
    .C(_2360_));
 sg13g2_a21oi_1 _3320_ (.A1(_2356_),
    .A2(_2360_),
    .Y(_2362_),
    .B1(_2354_));
 sg13g2_a21oi_1 _3321_ (.A1(_2303_),
    .A2(_2305_),
    .Y(_2363_),
    .B1(_2310_));
 sg13g2_a21oi_1 _3322_ (.A1(_2303_),
    .A2(_2305_),
    .Y(_2364_),
    .B1(_2311_));
 sg13g2_nor3_1 _3323_ (.A(_2302_),
    .B(_2304_),
    .C(_2310_),
    .Y(_2365_));
 sg13g2_nor3_1 _3324_ (.A(_2312_),
    .B(_2362_),
    .C(_2363_),
    .Y(_2366_));
 sg13g2_o21ai_1 _3325_ (.B1(_2358_),
    .Y(_2367_),
    .A1(_1460_),
    .A2(_2359_));
 sg13g2_inv_1 _3326_ (.Y(_2368_),
    .A(_2367_));
 sg13g2_nor4_1 _3327_ (.A(_2354_),
    .B(_2361_),
    .C(_2364_),
    .D(_2365_),
    .Y(_2369_));
 sg13g2_nor3_1 _3328_ (.A(_2366_),
    .B(_2368_),
    .C(_2369_),
    .Y(_2370_));
 sg13g2_nor2_1 _3329_ (.A(_2366_),
    .B(_2370_),
    .Y(_2371_));
 sg13g2_xnor2_1 _3330_ (.Y(_2372_),
    .A(_2316_),
    .B(_2317_));
 sg13g2_nand2_1 _3331_ (.Y(_2373_),
    .A(_2371_),
    .B(_2372_));
 sg13g2_o21ai_1 _3332_ (.B1(_2368_),
    .Y(_2374_),
    .A1(_2366_),
    .A2(_2369_));
 sg13g2_nand2b_1 _3333_ (.Y(_2375_),
    .B(_2374_),
    .A_N(_2370_));
 sg13g2_nand2_2 _3334_ (.Y(_2376_),
    .A(net652),
    .B(net512));
 sg13g2_nor2_2 _3335_ (.A(_2252_),
    .B(_2376_),
    .Y(_2377_));
 sg13g2_a22oi_1 _3336_ (.Y(_2378_),
    .B1(net509),
    .B2(net512),
    .A2(net510),
    .A1(net652));
 sg13g2_nor2_1 _3337_ (.A(_2377_),
    .B(_2378_),
    .Y(_2379_));
 sg13g2_nor2_1 _3338_ (.A(net512),
    .B(_2254_),
    .Y(_2380_));
 sg13g2_a21oi_1 _3339_ (.A1(_2252_),
    .A2(_2380_),
    .Y(_2381_),
    .B1(_2324_));
 sg13g2_nand2_1 _3340_ (.Y(_2382_),
    .A(_2266_),
    .B(_2341_));
 sg13g2_nand2_1 _3341_ (.Y(_2383_),
    .A(_2332_),
    .B(_2382_));
 sg13g2_nand3_1 _3342_ (.B(_2377_),
    .C(_2382_),
    .A(_2332_),
    .Y(_2384_));
 sg13g2_xor2_1 _3343_ (.B(_2383_),
    .A(_2377_),
    .X(_2385_));
 sg13g2_xnor2_1 _3344_ (.Y(_2386_),
    .A(_2379_),
    .B(_2381_));
 sg13g2_nor2_1 _3345_ (.A(_2385_),
    .B(_2386_),
    .Y(_2387_));
 sg13g2_a21oi_1 _3346_ (.A1(_2379_),
    .A2(_2381_),
    .Y(_2388_),
    .B1(_2387_));
 sg13g2_xor2_1 _3347_ (.B(_2336_),
    .A(_2328_),
    .X(_2389_));
 sg13g2_nor2b_1 _3348_ (.A(_2388_),
    .B_N(_2389_),
    .Y(_2390_));
 sg13g2_xnor2_1 _3349_ (.Y(_2391_),
    .A(_2388_),
    .B(_2389_));
 sg13g2_xor2_1 _3350_ (.B(_2342_),
    .A(_2341_),
    .X(_2392_));
 sg13g2_nand2_1 _3351_ (.Y(_2393_),
    .A(_2096_),
    .B(_2392_));
 sg13g2_xor2_1 _3352_ (.B(_2345_),
    .A(_2257_),
    .X(_2394_));
 sg13g2_nor2b_1 _3353_ (.A(_2384_),
    .B_N(_2394_),
    .Y(_2395_));
 sg13g2_xnor2_1 _3354_ (.Y(_2396_),
    .A(_2384_),
    .B(_2394_));
 sg13g2_nor2b_1 _3355_ (.A(_2393_),
    .B_N(_2396_),
    .Y(_2397_));
 sg13g2_xnor2_1 _3356_ (.Y(_2398_),
    .A(_2393_),
    .B(_2396_));
 sg13g2_a21oi_1 _3357_ (.A1(_2391_),
    .A2(_2398_),
    .Y(_2399_),
    .B1(_2390_));
 sg13g2_xor2_1 _3358_ (.B(_2351_),
    .A(_2340_),
    .X(_2400_));
 sg13g2_nor2b_1 _3359_ (.A(_2399_),
    .B_N(_2400_),
    .Y(_2401_));
 sg13g2_nor2_1 _3360_ (.A(_2395_),
    .B(_2397_),
    .Y(_2402_));
 sg13g2_nor2_1 _3361_ (.A(_0846_),
    .B(_2402_),
    .Y(_2403_));
 sg13g2_xnor2_1 _3362_ (.Y(_2404_),
    .A(_0835_),
    .B(_2402_));
 sg13g2_xnor2_1 _3363_ (.Y(_2405_),
    .A(_2399_),
    .B(_2400_));
 sg13g2_a21oi_1 _3364_ (.A1(_2404_),
    .A2(_2405_),
    .Y(_2406_),
    .B1(_2401_));
 sg13g2_a21oi_1 _3365_ (.A1(_2355_),
    .A2(_2356_),
    .Y(_2407_),
    .B1(_2360_));
 sg13g2_nor3_1 _3366_ (.A(_2361_),
    .B(_2406_),
    .C(_2407_),
    .Y(_2408_));
 sg13g2_or3_1 _3367_ (.A(_2361_),
    .B(_2406_),
    .C(_2407_),
    .X(_2409_));
 sg13g2_o21ai_1 _3368_ (.B1(_2406_),
    .Y(_2410_),
    .A1(_2361_),
    .A2(_2407_));
 sg13g2_nand3_1 _3369_ (.B(_2409_),
    .C(_2410_),
    .A(_2403_),
    .Y(_2411_));
 sg13g2_a21oi_1 _3370_ (.A1(_2403_),
    .A2(_2410_),
    .Y(_2412_),
    .B1(_2408_));
 sg13g2_a21o_1 _3371_ (.A2(_2410_),
    .A1(_2403_),
    .B1(_2408_),
    .X(_2413_));
 sg13g2_nand3b_1 _3372_ (.B(_2374_),
    .C(_2413_),
    .Y(_2414_),
    .A_N(_2370_));
 sg13g2_a21o_1 _3373_ (.A2(_2410_),
    .A1(_2409_),
    .B1(_2403_),
    .X(_2415_));
 sg13g2_nor3_1 _3374_ (.A(net509),
    .B(_2331_),
    .C(_2376_),
    .Y(_2416_));
 sg13g2_xor2_1 _3375_ (.B(_2386_),
    .A(_2385_),
    .X(_2417_));
 sg13g2_nand2_1 _3376_ (.Y(_2418_),
    .A(_2416_),
    .B(_2417_));
 sg13g2_xor2_1 _3377_ (.B(_2417_),
    .A(_2416_),
    .X(_2419_));
 sg13g2_xnor2_1 _3378_ (.Y(_2420_),
    .A(_2613_),
    .B(net537));
 sg13g2_xnor2_1 _3379_ (.Y(_2421_),
    .A(net596),
    .B(net536));
 sg13g2_nor2_2 _3380_ (.A(_2635_),
    .B(_2420_),
    .Y(_2422_));
 sg13g2_nand2_1 _3381_ (.Y(_2423_),
    .A(net497),
    .B(_2422_));
 sg13g2_or3_1 _3382_ (.A(_1032_),
    .B(_2331_),
    .C(_2376_),
    .X(_2424_));
 sg13g2_xnor2_1 _3383_ (.Y(_2425_),
    .A(_2097_),
    .B(_2392_));
 sg13g2_nor2b_1 _3384_ (.A(_2424_),
    .B_N(_2425_),
    .Y(_2426_));
 sg13g2_xor2_1 _3385_ (.B(_2425_),
    .A(_2424_),
    .X(_2427_));
 sg13g2_nor2_1 _3386_ (.A(_2423_),
    .B(_2427_),
    .Y(_2428_));
 sg13g2_xor2_1 _3387_ (.B(_2427_),
    .A(_2423_),
    .X(_2429_));
 sg13g2_nand2_1 _3388_ (.Y(_2430_),
    .A(_2419_),
    .B(_2429_));
 sg13g2_nand2_1 _3389_ (.Y(_2431_),
    .A(_2418_),
    .B(_2430_));
 sg13g2_xnor2_1 _3390_ (.Y(_2432_),
    .A(_2391_),
    .B(_2398_));
 sg13g2_nor2b_1 _3391_ (.A(_2432_),
    .B_N(_2431_),
    .Y(_2433_));
 sg13g2_o21ai_1 _3392_ (.B1(_2256_),
    .Y(_2434_),
    .A1(_2426_),
    .A2(_2428_));
 sg13g2_or3_1 _3393_ (.A(_2256_),
    .B(_2426_),
    .C(_2428_),
    .X(_2435_));
 sg13g2_and2_1 _3394_ (.A(_2434_),
    .B(_2435_),
    .X(_2436_));
 sg13g2_xnor2_1 _3395_ (.Y(_2437_),
    .A(_2431_),
    .B(_2432_));
 sg13g2_a21oi_1 _3396_ (.A1(_2436_),
    .A2(_2437_),
    .Y(_2438_),
    .B1(_2433_));
 sg13g2_xnor2_1 _3397_ (.Y(_2439_),
    .A(_2404_),
    .B(_2405_));
 sg13g2_or2_1 _3398_ (.X(_2440_),
    .B(_2439_),
    .A(_2438_));
 sg13g2_and2_1 _3399_ (.A(_2438_),
    .B(_2439_),
    .X(_2441_));
 sg13g2_xor2_1 _3400_ (.B(_2439_),
    .A(_2438_),
    .X(_2442_));
 sg13g2_o21ai_1 _3401_ (.B1(_2440_),
    .Y(_2443_),
    .A1(_2434_),
    .A2(_2441_));
 sg13g2_nand3_1 _3402_ (.B(_2415_),
    .C(_2443_),
    .A(_2411_),
    .Y(_2444_));
 sg13g2_xnor2_1 _3403_ (.Y(_2445_),
    .A(_2436_),
    .B(_2437_));
 sg13g2_nor2_2 _3404_ (.A(net561),
    .B(_2613_),
    .Y(_2446_));
 sg13g2_nand2_2 _3405_ (.Y(_2447_),
    .A(net592),
    .B(net595));
 sg13g2_nor2_2 _3406_ (.A(_1262_),
    .B(_2446_),
    .Y(_2448_));
 sg13g2_nand2_2 _3407_ (.Y(_2449_),
    .A(_1273_),
    .B(_2447_));
 sg13g2_nor2_1 _3408_ (.A(_1875_),
    .B(_2449_),
    .Y(_2450_));
 sg13g2_nor2_1 _3409_ (.A(_2419_),
    .B(_2429_),
    .Y(_2451_));
 sg13g2_xor2_1 _3410_ (.B(_2376_),
    .A(_2331_),
    .X(_2452_));
 sg13g2_nand3_1 _3411_ (.B(net509),
    .C(_2452_),
    .A(net653),
    .Y(_2453_));
 sg13g2_mux2_1 _3412_ (.A0(net507),
    .A1(_1875_),
    .S(_2449_),
    .X(_2454_));
 sg13g2_a21oi_1 _3413_ (.A1(net653),
    .A2(net509),
    .Y(_2455_),
    .B1(_2452_));
 sg13g2_o21ai_1 _3414_ (.B1(_2453_),
    .Y(_2456_),
    .A1(_2454_),
    .A2(_2455_));
 sg13g2_xnor2_1 _3415_ (.Y(_2457_),
    .A(_2255_),
    .B(_2450_));
 sg13g2_nor2_1 _3416_ (.A(_2456_),
    .B(_2457_),
    .Y(_2458_));
 sg13g2_nor2_1 _3417_ (.A(_2451_),
    .B(_2458_),
    .Y(_2459_));
 sg13g2_a22oi_1 _3418_ (.Y(_2460_),
    .B1(_2459_),
    .B2(_2430_),
    .A2(_2457_),
    .A1(_2456_));
 sg13g2_xnor2_1 _3419_ (.Y(_2461_),
    .A(_2445_),
    .B(_2460_));
 sg13g2_nor4_1 _3420_ (.A(_1875_),
    .B(_2255_),
    .C(_2449_),
    .D(_2461_),
    .Y(_2462_));
 sg13g2_nor2_1 _3421_ (.A(_2445_),
    .B(_2460_),
    .Y(_2463_));
 sg13g2_xnor2_1 _3422_ (.Y(_2464_),
    .A(_2434_),
    .B(_2442_));
 sg13g2_o21ai_1 _3423_ (.B1(_2464_),
    .Y(_2465_),
    .A1(_2462_),
    .A2(_2463_));
 sg13g2_a21oi_1 _3424_ (.A1(_2411_),
    .A2(_2415_),
    .Y(_2466_),
    .B1(_2443_));
 sg13g2_a221oi_1 _3425_ (.B2(_2465_),
    .C1(_2466_),
    .B1(_2444_),
    .A1(_2375_),
    .Y(_2467_),
    .A2(_2412_));
 sg13g2_xor2_1 _3426_ (.B(_2372_),
    .A(_2371_),
    .X(_2468_));
 sg13g2_o21ai_1 _3427_ (.B1(_2414_),
    .Y(_2469_),
    .A1(_2371_),
    .A2(_2372_));
 sg13g2_a22oi_1 _3428_ (.Y(_2470_),
    .B1(_2469_),
    .B2(_2373_),
    .A2(_2468_),
    .A1(_2467_));
 sg13g2_and2_1 _3429_ (.A(_2251_),
    .B(_2318_),
    .X(_2471_));
 sg13g2_or2_1 _3430_ (.X(_2472_),
    .B(_2471_),
    .A(_2249_));
 sg13g2_nor2_1 _3431_ (.A(_2249_),
    .B(_2321_),
    .Y(_2473_));
 sg13g2_o21ai_1 _3432_ (.B1(_2322_),
    .Y(_2474_),
    .A1(_2470_),
    .A2(_2472_));
 sg13g2_a21oi_1 _3433_ (.A1(_2217_),
    .A2(_2218_),
    .Y(_2475_),
    .B1(_2220_));
 sg13g2_a21o_1 _3434_ (.A2(_2243_),
    .A1(_2221_),
    .B1(_2242_),
    .X(_2476_));
 sg13g2_and2_1 _3435_ (.A(_2064_),
    .B(_2223_),
    .X(_2477_));
 sg13g2_xnor2_1 _3436_ (.Y(_2478_),
    .A(_2064_),
    .B(_2223_));
 sg13g2_inv_1 _3437_ (.Y(_2479_),
    .A(_2478_));
 sg13g2_a21oi_1 _3438_ (.A1(_2224_),
    .A2(_2240_),
    .Y(_2480_),
    .B1(_2239_));
 sg13g2_o21ai_1 _3439_ (.B1(_2236_),
    .Y(_2481_),
    .A1(_2231_),
    .A2(_2237_));
 sg13g2_o21ai_1 _3440_ (.B1(_2233_),
    .Y(_2482_),
    .A1(_2098_),
    .A2(_2234_));
 sg13g2_o21ai_1 _3441_ (.B1(net462),
    .Y(_2483_),
    .A1(_2027_),
    .A2(_2228_));
 sg13g2_xor2_1 _3442_ (.B(_2483_),
    .A(_2482_),
    .X(_2484_));
 sg13g2_inv_1 _3443_ (.Y(_2485_),
    .A(_2484_));
 sg13g2_nand2_1 _3444_ (.Y(_2486_),
    .A(_2481_),
    .B(_2485_));
 sg13g2_xnor2_1 _3445_ (.Y(_2487_),
    .A(_2481_),
    .B(_2484_));
 sg13g2_nor2_1 _3446_ (.A(_0978_),
    .B(_2230_),
    .Y(_2488_));
 sg13g2_xnor2_1 _3447_ (.Y(_2489_),
    .A(_0978_),
    .B(_2230_));
 sg13g2_inv_1 _3448_ (.Y(_2490_),
    .A(_2489_));
 sg13g2_nand2_1 _3449_ (.Y(_2491_),
    .A(_2487_),
    .B(_2490_));
 sg13g2_xnor2_1 _3450_ (.Y(_2492_),
    .A(_2487_),
    .B(_2490_));
 sg13g2_nor2_1 _3451_ (.A(_2480_),
    .B(_2492_),
    .Y(_2493_));
 sg13g2_xor2_1 _3452_ (.B(_2492_),
    .A(_2480_),
    .X(_2494_));
 sg13g2_xnor2_1 _3453_ (.Y(_2495_),
    .A(_2478_),
    .B(_2494_));
 sg13g2_nand2_1 _3454_ (.Y(_2496_),
    .A(_2476_),
    .B(_2495_));
 sg13g2_xor2_1 _3455_ (.B(_2495_),
    .A(_2476_),
    .X(_2497_));
 sg13g2_nand2b_1 _3456_ (.Y(_2498_),
    .B(_2497_),
    .A_N(_2475_));
 sg13g2_xor2_1 _3457_ (.B(_2497_),
    .A(_2475_),
    .X(_2499_));
 sg13g2_a21oi_1 _3458_ (.A1(_2215_),
    .A2(_2247_),
    .Y(_2500_),
    .B1(_2245_));
 sg13g2_nor2_1 _3459_ (.A(_2499_),
    .B(_2500_),
    .Y(_2501_));
 sg13g2_xor2_1 _3460_ (.B(_2500_),
    .A(_2499_),
    .X(_2502_));
 sg13g2_xnor2_1 _3461_ (.Y(_2503_),
    .A(_2474_),
    .B(_2502_));
 sg13g2_a21oi_1 _3462_ (.A1(_2479_),
    .A2(_2494_),
    .Y(_2504_),
    .B1(_2493_));
 sg13g2_nand2_1 _3463_ (.Y(_2505_),
    .A(_1065_),
    .B(_1799_));
 sg13g2_nor3_1 _3464_ (.A(_0978_),
    .B(_2230_),
    .C(_2505_),
    .Y(_2506_));
 sg13g2_xnor2_1 _3465_ (.Y(_2507_),
    .A(_2488_),
    .B(_2505_));
 sg13g2_nand2_1 _3466_ (.Y(_2508_),
    .A(net462),
    .B(_2482_));
 sg13g2_nor2_1 _3467_ (.A(_2228_),
    .B(_2508_),
    .Y(_2509_));
 sg13g2_xnor2_1 _3468_ (.Y(_2510_),
    .A(_2228_),
    .B(_2508_));
 sg13g2_a21oi_1 _3469_ (.A1(_2486_),
    .A2(_2491_),
    .Y(_2511_),
    .B1(_2510_));
 sg13g2_nand3_1 _3470_ (.B(_2491_),
    .C(_2510_),
    .A(_2486_),
    .Y(_2512_));
 sg13g2_nor2b_1 _3471_ (.A(_2511_),
    .B_N(_2512_),
    .Y(_2513_));
 sg13g2_xnor2_1 _3472_ (.Y(_2514_),
    .A(_2507_),
    .B(_2513_));
 sg13g2_nor2_1 _3473_ (.A(_2504_),
    .B(_2514_),
    .Y(_2515_));
 sg13g2_xor2_1 _3474_ (.B(_2514_),
    .A(_2504_),
    .X(_2516_));
 sg13g2_xnor2_1 _3475_ (.Y(_2517_),
    .A(_2477_),
    .B(_2516_));
 sg13g2_nand3_1 _3476_ (.B(_2498_),
    .C(_2517_),
    .A(_2496_),
    .Y(_2518_));
 sg13g2_inv_1 _3477_ (.Y(_2519_),
    .A(_2518_));
 sg13g2_a21o_1 _3478_ (.A2(_2498_),
    .A1(_2496_),
    .B1(_2517_),
    .X(_2520_));
 sg13g2_and2_1 _3479_ (.A(_2518_),
    .B(_2520_),
    .X(_2521_));
 sg13g2_a21oi_1 _3480_ (.A1(_2474_),
    .A2(_2502_),
    .Y(_2522_),
    .B1(_2501_));
 sg13g2_xor2_1 _3481_ (.B(_2522_),
    .A(_2521_),
    .X(_2523_));
 sg13g2_xnor2_1 _3482_ (.Y(_2524_),
    .A(_2521_),
    .B(_2522_));
 sg13g2_and2_1 _3483_ (.A(_2503_),
    .B(_2523_),
    .X(_2525_));
 sg13g2_nand2b_1 _3484_ (.Y(_2526_),
    .B(_2520_),
    .A_N(_2501_));
 sg13g2_a21oi_1 _3485_ (.A1(_2474_),
    .A2(_2502_),
    .Y(_2527_),
    .B1(_2526_));
 sg13g2_a21o_1 _3486_ (.A2(_2502_),
    .A1(_2474_),
    .B1(_2526_),
    .X(_2528_));
 sg13g2_a21oi_1 _3487_ (.A1(_2477_),
    .A2(_2516_),
    .Y(_2529_),
    .B1(_2515_));
 sg13g2_xor2_1 _3488_ (.B(_2511_),
    .A(_2506_),
    .X(_2530_));
 sg13g2_a21oi_1 _3489_ (.A1(_2507_),
    .A2(_2513_),
    .Y(_2531_),
    .B1(_2530_));
 sg13g2_nor2_1 _3490_ (.A(net463),
    .B(_1581_),
    .Y(_2532_));
 sg13g2_inv_1 _3491_ (.Y(_2533_),
    .A(_2532_));
 sg13g2_nand2_1 _3492_ (.Y(_2534_),
    .A(_0978_),
    .B(net461));
 sg13g2_xnor2_1 _3493_ (.Y(_2535_),
    .A(_2532_),
    .B(_2534_));
 sg13g2_xnor2_1 _3494_ (.Y(_2536_),
    .A(_2509_),
    .B(_2535_));
 sg13g2_xnor2_1 _3495_ (.Y(_2537_),
    .A(_2531_),
    .B(_2536_));
 sg13g2_xor2_1 _3496_ (.B(_2537_),
    .A(_2529_),
    .X(_2538_));
 sg13g2_inv_1 _3497_ (.Y(_2539_),
    .A(_2538_));
 sg13g2_nand3_1 _3498_ (.B(_2528_),
    .C(_2538_),
    .A(_2518_),
    .Y(_2540_));
 sg13g2_o21ai_1 _3499_ (.B1(_2539_),
    .Y(_2541_),
    .A1(_2519_),
    .A2(_2527_));
 sg13g2_nand3_1 _3500_ (.B(_2528_),
    .C(_2539_),
    .A(_2518_),
    .Y(_2542_));
 sg13g2_o21ai_1 _3501_ (.B1(_2538_),
    .Y(_2543_),
    .A1(_2519_),
    .A2(_2527_));
 sg13g2_nand2_2 _3502_ (.Y(_2544_),
    .A(_2542_),
    .B(_2543_));
 sg13g2_a22oi_1 _3503_ (.Y(_2545_),
    .B1(_2542_),
    .B2(_2543_),
    .A2(_2523_),
    .A1(_2503_));
 sg13g2_o21ai_1 _3504_ (.B1(_2320_),
    .Y(_2546_),
    .A1(_2470_),
    .A2(_2471_));
 sg13g2_xnor2_1 _3505_ (.Y(_2547_),
    .A(_2473_),
    .B(_2546_));
 sg13g2_nand2_1 _3506_ (.Y(_2548_),
    .A(_2503_),
    .B(_2547_));
 sg13g2_a22oi_1 _3507_ (.Y(_2549_),
    .B1(_2548_),
    .B2(_2524_),
    .A2(_2541_),
    .A1(_2540_));
 sg13g2_nand2_1 _3508_ (.Y(_2550_),
    .A(_2227_),
    .B(_2228_));
 sg13g2_nor2_1 _3509_ (.A(_2112_),
    .B(_2550_),
    .Y(_2551_));
 sg13g2_nor2_2 _3510_ (.A(net556),
    .B(net555),
    .Y(_2552_));
 sg13g2_nand2_2 _3511_ (.Y(_2553_),
    .A(net625),
    .B(net620));
 sg13g2_nand3_1 _3512_ (.B(_0923_),
    .C(_2552_),
    .A(net612),
    .Y(_2554_));
 sg13g2_nand2_2 _3513_ (.Y(_2555_),
    .A(_2712_),
    .B(net553));
 sg13g2_and2_1 _3514_ (.A(net634),
    .B(net629),
    .X(_2556_));
 sg13g2_nand2_2 _3515_ (.Y(_2557_),
    .A(net632),
    .B(net631));
 sg13g2_nor2_1 _3516_ (.A(_2555_),
    .B(_2556_),
    .Y(_2559_));
 sg13g2_nor3_1 _3517_ (.A(net607),
    .B(_0604_),
    .C(_2559_),
    .Y(_2560_));
 sg13g2_nand3_1 _3518_ (.B(_2554_),
    .C(_2560_),
    .A(_2551_),
    .Y(_2561_));
 sg13g2_nor3_1 _3519_ (.A(_2545_),
    .B(_2549_),
    .C(_2561_),
    .Y(_2562_));
 sg13g2_or3_1 _3520_ (.A(_2545_),
    .B(_2549_),
    .C(_2561_),
    .X(_2563_));
 sg13g2_nor2b_2 _3521_ (.A(net550),
    .B_N(_0076_),
    .Y(_2564_));
 sg13g2_nor2b_2 _3522_ (.A(_0087_),
    .B_N(_2564_),
    .Y(_2565_));
 sg13g2_nand2b_2 _3523_ (.Y(_2566_),
    .B(_2564_),
    .A_N(_0087_));
 sg13g2_nor2b_2 _3524_ (.A(_0142_),
    .B_N(_0131_),
    .Y(_2567_));
 sg13g2_nand2_2 _3525_ (.Y(_2568_),
    .A(_0296_),
    .B(_2567_));
 sg13g2_nor2_2 _3526_ (.A(net496),
    .B(_2568_),
    .Y(_2570_));
 sg13g2_and2_1 _3527_ (.A(_2563_),
    .B(_2570_),
    .X(_2571_));
 sg13g2_nor2_2 _3528_ (.A(net577),
    .B(net583),
    .Y(_2572_));
 sg13g2_o21ai_1 _3529_ (.B1(net572),
    .Y(_2573_),
    .A1(net579),
    .A2(net582));
 sg13g2_and2_1 _3530_ (.A(net562),
    .B(_2573_),
    .X(_2574_));
 sg13g2_nand2_1 _3531_ (.Y(_2575_),
    .A(net564),
    .B(_2573_));
 sg13g2_and2_1 _3532_ (.A(_0439_),
    .B(_2567_),
    .X(_2576_));
 sg13g2_nand2_2 _3533_ (.Y(_2577_),
    .A(_0439_),
    .B(_2567_));
 sg13g2_nand2_2 _3534_ (.Y(_2578_),
    .A(_2565_),
    .B(_2576_));
 sg13g2_nor2_1 _3535_ (.A(net526),
    .B(_2578_),
    .Y(_2579_));
 sg13g2_nor2_1 _3536_ (.A(_2635_),
    .B(net559),
    .Y(_2581_));
 sg13g2_nand2_2 _3537_ (.Y(_2582_),
    .A(net603),
    .B(net653));
 sg13g2_nor2_2 _3538_ (.A(net604),
    .B(net652),
    .Y(_2583_));
 sg13g2_nand2_2 _3539_ (.Y(_2584_),
    .A(_2635_),
    .B(net559));
 sg13g2_nor2_2 _3540_ (.A(_2581_),
    .B(_2583_),
    .Y(_2585_));
 sg13g2_nand2_1 _3541_ (.Y(_2586_),
    .A(_2582_),
    .B(_2584_));
 sg13g2_nor2_1 _3542_ (.A(net573),
    .B(net578),
    .Y(_2587_));
 sg13g2_nor2_1 _3543_ (.A(net563),
    .B(_2587_),
    .Y(_2588_));
 sg13g2_o21ai_1 _3544_ (.B1(net570),
    .Y(_2589_),
    .A1(net576),
    .A2(net581));
 sg13g2_nand2_2 _3545_ (.Y(_2590_),
    .A(net484),
    .B(net523));
 sg13g2_a21oi_1 _3546_ (.A1(net527),
    .A2(_2590_),
    .Y(_2592_),
    .B1(_2578_));
 sg13g2_a21oi_1 _3547_ (.A1(_2563_),
    .A2(_2570_),
    .Y(_2593_),
    .B1(_2592_));
 sg13g2_nand2_2 _3548_ (.Y(_2594_),
    .A(net618),
    .B(net612));
 sg13g2_nor2_1 _3549_ (.A(net618),
    .B(net606),
    .Y(_2595_));
 sg13g2_a21oi_2 _3550_ (.B1(net608),
    .Y(_2596_),
    .A2(_2552_),
    .A1(net611));
 sg13g2_o21ai_1 _3551_ (.B1(_2596_),
    .Y(_2597_),
    .A1(net612),
    .A2(_2552_));
 sg13g2_nand2b_1 _3552_ (.Y(_2598_),
    .B(_1581_),
    .A_N(_2597_));
 sg13g2_a221oi_1 _3553_ (.B2(_2524_),
    .C1(_2598_),
    .B1(_2548_),
    .A1(_2540_),
    .Y(_2599_),
    .A2(_2541_));
 sg13g2_nand3b_1 _3554_ (.B(_1581_),
    .C(_2549_),
    .Y(_2600_),
    .A_N(_2597_));
 sg13g2_a21o_2 _3555_ (.A2(_2599_),
    .A1(_2525_),
    .B1(_0241_),
    .X(_2601_));
 sg13g2_nor2_2 _3556_ (.A(net566),
    .B(net574),
    .Y(_2603_));
 sg13g2_or2_1 _3557_ (.X(_2604_),
    .B(net574),
    .A(net568));
 sg13g2_nand2_2 _3558_ (.Y(_2605_),
    .A(_2569_),
    .B(_0527_));
 sg13g2_nor2_2 _3559_ (.A(_0516_),
    .B(_2604_),
    .Y(_2606_));
 sg13g2_nand2_2 _3560_ (.Y(_2607_),
    .A(_0527_),
    .B(net541));
 sg13g2_nor2_1 _3561_ (.A(net490),
    .B(net522),
    .Y(_2608_));
 sg13g2_o21ai_1 _3562_ (.B1(_1098_),
    .Y(_2609_),
    .A1(_1152_),
    .A2(_2447_));
 sg13g2_nand2_1 _3563_ (.Y(_2610_),
    .A(net549),
    .B(_2609_));
 sg13g2_or2_1 _3564_ (.X(_2611_),
    .B(_2609_),
    .A(net491));
 sg13g2_a21oi_1 _3565_ (.A1(_2610_),
    .A2(_2611_),
    .Y(_2612_),
    .B1(_2606_));
 sg13g2_nand2_2 _3566_ (.Y(_2614_),
    .A(net494),
    .B(_2606_));
 sg13g2_nor2b_1 _3567_ (.A(_2612_),
    .B_N(_2614_),
    .Y(_2615_));
 sg13g2_a21o_1 _3568_ (.A2(_2615_),
    .A1(_2600_),
    .B1(_2601_),
    .X(_2616_));
 sg13g2_and4_1 _3569_ (.A(_2105_),
    .B(_2195_),
    .C(_2505_),
    .D(_2551_),
    .X(_2617_));
 sg13g2_and3_1 _3570_ (.X(_2618_),
    .A(_2503_),
    .B(_2523_),
    .C(_2617_));
 sg13g2_and2_1 _3571_ (.A(_2544_),
    .B(_2618_),
    .X(_2619_));
 sg13g2_nor2_1 _3572_ (.A(net555),
    .B(net612),
    .Y(_2620_));
 sg13g2_or2_1 _3573_ (.X(_2621_),
    .B(_1799_),
    .A(_1570_));
 sg13g2_nor2_1 _3574_ (.A(_2544_),
    .B(_2621_),
    .Y(_2622_));
 sg13g2_o21ai_1 _3575_ (.B1(_2620_),
    .Y(_2623_),
    .A1(_2544_),
    .A2(_2621_));
 sg13g2_and2_1 _3576_ (.A(_0131_),
    .B(_0142_),
    .X(_2625_));
 sg13g2_nand2_2 _3577_ (.Y(_2626_),
    .A(_0439_),
    .B(_2625_));
 sg13g2_and2_1 _3578_ (.A(_0087_),
    .B(_2564_),
    .X(_2627_));
 sg13g2_nand2_2 _3579_ (.Y(_2628_),
    .A(_0087_),
    .B(_2564_));
 sg13g2_nor2_2 _3580_ (.A(_2626_),
    .B(net478),
    .Y(_2629_));
 sg13g2_nor3_1 _3581_ (.A(net608),
    .B(_2626_),
    .C(net478),
    .Y(_2630_));
 sg13g2_o21ai_1 _3582_ (.B1(_2630_),
    .Y(_2631_),
    .A1(_2619_),
    .A2(_2623_));
 sg13g2_nor2_1 _3583_ (.A(_2042_),
    .B(_2155_),
    .Y(_2632_));
 sg13g2_a21oi_1 _3584_ (.A1(_2027_),
    .A2(_2042_),
    .Y(_2633_),
    .B1(_2049_));
 sg13g2_nand2b_2 _3585_ (.Y(_2634_),
    .B(_2633_),
    .A_N(_2632_));
 sg13g2_nand2_2 _3586_ (.Y(_2636_),
    .A(net631),
    .B(net625));
 sg13g2_inv_1 _3587_ (.Y(_2637_),
    .A(_2636_));
 sg13g2_nor3_2 _3588_ (.A(net620),
    .B(net615),
    .C(net610),
    .Y(_2638_));
 sg13g2_or3_1 _3589_ (.A(net620),
    .B(net615),
    .C(net610),
    .X(_2639_));
 sg13g2_and2_1 _3590_ (.A(_2636_),
    .B(_2638_),
    .X(_2640_));
 sg13g2_and2_1 _3591_ (.A(net644),
    .B(net639),
    .X(_2641_));
 sg13g2_nand2_1 _3592_ (.Y(_2642_),
    .A(net645),
    .B(net639));
 sg13g2_a21oi_2 _3593_ (.B1(net636),
    .Y(_2643_),
    .A2(net639),
    .A1(net643));
 sg13g2_o21ai_1 _3594_ (.B1(net625),
    .Y(_2644_),
    .A1(_0945_),
    .A2(_2641_));
 sg13g2_nand2_2 _3595_ (.Y(_2645_),
    .A(_2640_),
    .B(_2644_));
 sg13g2_nand2_2 _3596_ (.Y(_2647_),
    .A(net649),
    .B(net639));
 sg13g2_and3_1 _3597_ (.X(_2648_),
    .A(net649),
    .B(net643),
    .C(net639));
 sg13g2_nand3_1 _3598_ (.B(net643),
    .C(net639),
    .A(net649),
    .Y(_2649_));
 sg13g2_nand2_1 _3599_ (.Y(_2650_),
    .A(net547),
    .B(_2649_));
 sg13g2_and3_1 _3600_ (.X(_2651_),
    .A(_2640_),
    .B(_2644_),
    .C(_2650_));
 sg13g2_nand3_1 _3601_ (.B(_2644_),
    .C(_2650_),
    .A(_2640_),
    .Y(_2652_));
 sg13g2_nor3_1 _3602_ (.A(_0945_),
    .B(_2640_),
    .C(_2641_),
    .Y(_2653_));
 sg13g2_o21ai_1 _3603_ (.B1(net631),
    .Y(_2654_),
    .A1(_2651_),
    .A2(_2653_));
 sg13g2_or3_1 _3604_ (.A(net631),
    .B(_2651_),
    .C(_2653_),
    .X(_2655_));
 sg13g2_and2_1 _3605_ (.A(_2654_),
    .B(_2655_),
    .X(_2656_));
 sg13g2_inv_1 _3606_ (.Y(_2658_),
    .A(_2656_));
 sg13g2_and3_1 _3607_ (.X(_2659_),
    .A(net648),
    .B(_2654_),
    .C(_2655_));
 sg13g2_a21o_2 _3608_ (.A2(_2659_),
    .A1(_2271_),
    .B1(_2268_),
    .X(_2660_));
 sg13g2_xnor2_1 _3609_ (.Y(_2661_),
    .A(_2042_),
    .B(_2049_));
 sg13g2_nor2b_1 _3610_ (.A(_2661_),
    .B_N(_2660_),
    .Y(_2662_));
 sg13g2_xnor2_1 _3611_ (.Y(_2663_),
    .A(net632),
    .B(_2643_));
 sg13g2_a21o_1 _3612_ (.A2(_2644_),
    .A1(_2640_),
    .B1(_2663_),
    .X(_2664_));
 sg13g2_a21oi_1 _3613_ (.A1(net558),
    .A2(_2649_),
    .Y(_2665_),
    .B1(net557));
 sg13g2_o21ai_1 _3614_ (.B1(_2664_),
    .Y(_2666_),
    .A1(_2652_),
    .A2(_2665_));
 sg13g2_nor2_2 _3615_ (.A(net558),
    .B(_2690_),
    .Y(_2667_));
 sg13g2_nand3_1 _3616_ (.B(net636),
    .C(net640),
    .A(net644),
    .Y(_2669_));
 sg13g2_and4_1 _3617_ (.A(net649),
    .B(net643),
    .C(net636),
    .D(net640),
    .X(_2670_));
 sg13g2_or2_1 _3618_ (.X(_2671_),
    .B(_2669_),
    .A(net559));
 sg13g2_a21oi_1 _3619_ (.A1(net558),
    .A2(_2649_),
    .Y(_2672_),
    .B1(_2670_));
 sg13g2_o21ai_1 _3620_ (.B1(_2671_),
    .Y(_2673_),
    .A1(net636),
    .A2(_2648_));
 sg13g2_nand2b_2 _3621_ (.Y(_2674_),
    .B(_2669_),
    .A_N(_2643_));
 sg13g2_nor2_1 _3622_ (.A(_2645_),
    .B(_2673_),
    .Y(_2675_));
 sg13g2_mux2_1 _3623_ (.A0(_2672_),
    .A1(_2674_),
    .S(_2645_),
    .X(_2676_));
 sg13g2_a21oi_1 _3624_ (.A1(_2645_),
    .A2(_2674_),
    .Y(_2677_),
    .B1(_2675_));
 sg13g2_a21oi_1 _3625_ (.A1(net649),
    .A2(net643),
    .Y(_2678_),
    .B1(net639));
 sg13g2_nor2_1 _3626_ (.A(_2648_),
    .B(_2678_),
    .Y(_2680_));
 sg13g2_or2_1 _3627_ (.X(_2681_),
    .B(_2678_),
    .A(_2648_));
 sg13g2_nor2_1 _3628_ (.A(_0692_),
    .B(_2641_),
    .Y(_2682_));
 sg13g2_nand2b_1 _3629_ (.Y(_2683_),
    .B(_2642_),
    .A_N(_0692_));
 sg13g2_mux2_1 _3630_ (.A0(_2681_),
    .A1(_2682_),
    .S(_2645_),
    .X(_2684_));
 sg13g2_nand2_2 _3631_ (.Y(_2685_),
    .A(_2666_),
    .B(_2684_));
 sg13g2_nand3_1 _3632_ (.B(net459),
    .C(_2684_),
    .A(_2666_),
    .Y(_2686_));
 sg13g2_xnor2_1 _3633_ (.Y(_2687_),
    .A(net459),
    .B(_2685_));
 sg13g2_xnor2_1 _3634_ (.Y(_2688_),
    .A(_2660_),
    .B(_2661_));
 sg13g2_a21oi_1 _3635_ (.A1(_2687_),
    .A2(_2688_),
    .Y(_2689_),
    .B1(_2662_));
 sg13g2_nor2_1 _3636_ (.A(_2634_),
    .B(_2689_),
    .Y(_2691_));
 sg13g2_xor2_1 _3637_ (.B(_2689_),
    .A(_2634_),
    .X(_2692_));
 sg13g2_nand2_2 _3638_ (.Y(_2693_),
    .A(_2656_),
    .B(_2684_));
 sg13g2_inv_1 _3639_ (.Y(_2694_),
    .A(_2693_));
 sg13g2_mux2_1 _3640_ (.A0(_1021_),
    .A1(_2668_),
    .S(_2645_),
    .X(_2695_));
 sg13g2_and2_1 _3641_ (.A(_2656_),
    .B(net458),
    .X(_2696_));
 sg13g2_nand2_2 _3642_ (.Y(_2697_),
    .A(_2656_),
    .B(_2666_));
 sg13g2_nand2_1 _3643_ (.Y(_2698_),
    .A(_2684_),
    .B(net458));
 sg13g2_nor2_1 _3644_ (.A(_2697_),
    .B(_2698_),
    .Y(_2699_));
 sg13g2_xnor2_1 _3645_ (.Y(_2700_),
    .A(_2685_),
    .B(_2696_));
 sg13g2_a21oi_1 _3646_ (.A1(_2043_),
    .A2(_2700_),
    .Y(_2702_),
    .B1(_2699_));
 sg13g2_nor2_1 _3647_ (.A(net460),
    .B(_2693_),
    .Y(_2703_));
 sg13g2_xor2_1 _3648_ (.B(_2693_),
    .A(net460),
    .X(_2704_));
 sg13g2_nor2b_1 _3649_ (.A(_2686_),
    .B_N(_2704_),
    .Y(_2705_));
 sg13g2_xnor2_1 _3650_ (.Y(_2706_),
    .A(_2686_),
    .B(_2704_));
 sg13g2_nor2b_1 _3651_ (.A(_2702_),
    .B_N(_2706_),
    .Y(_2707_));
 sg13g2_xnor2_1 _3652_ (.Y(_2708_),
    .A(_2702_),
    .B(_2706_));
 sg13g2_a21oi_1 _3653_ (.A1(_2692_),
    .A2(_2708_),
    .Y(_2709_),
    .B1(_2691_));
 sg13g2_nand2_1 _3654_ (.Y(_2710_),
    .A(_2666_),
    .B(net459));
 sg13g2_nor2_1 _3655_ (.A(_2142_),
    .B(_2710_),
    .Y(_2711_));
 sg13g2_nand2_1 _3656_ (.Y(_2713_),
    .A(_2142_),
    .B(_2710_));
 sg13g2_nand2b_1 _3657_ (.Y(_2714_),
    .B(_2713_),
    .A_N(_2711_));
 sg13g2_xor2_1 _3658_ (.B(_2714_),
    .A(_2703_),
    .X(_2715_));
 sg13g2_nor2_1 _3659_ (.A(_2677_),
    .B(_2697_),
    .Y(_2716_));
 sg13g2_nand2_1 _3660_ (.Y(_2717_),
    .A(_2656_),
    .B(_2676_));
 sg13g2_a21oi_1 _3661_ (.A1(_2656_),
    .A2(_2676_),
    .Y(_2718_),
    .B1(_2666_));
 sg13g2_or2_1 _3662_ (.X(_2719_),
    .B(_2718_),
    .A(_2716_));
 sg13g2_nor2b_1 _3663_ (.A(_2142_),
    .B_N(_2028_),
    .Y(_2720_));
 sg13g2_nor2_1 _3664_ (.A(_2142_),
    .B(_2719_),
    .Y(_2721_));
 sg13g2_xnor2_1 _3665_ (.Y(_2722_),
    .A(_2719_),
    .B(_2720_));
 sg13g2_nor2b_1 _3666_ (.A(_2715_),
    .B_N(_2722_),
    .Y(_2724_));
 sg13g2_xnor2_1 _3667_ (.Y(_2725_),
    .A(_2715_),
    .B(_2722_));
 sg13g2_inv_1 _3668_ (.Y(_2726_),
    .A(_2725_));
 sg13g2_nor2_1 _3669_ (.A(_2027_),
    .B(_2717_),
    .Y(_2727_));
 sg13g2_xnor2_1 _3670_ (.Y(_2728_),
    .A(net505),
    .B(_2717_));
 sg13g2_o21ai_1 _3671_ (.B1(_2728_),
    .Y(_2729_),
    .A1(_2705_),
    .A2(_2707_));
 sg13g2_or3_1 _3672_ (.A(_2705_),
    .B(_2707_),
    .C(_2728_),
    .X(_2730_));
 sg13g2_nand2_1 _3673_ (.Y(_2731_),
    .A(_2729_),
    .B(_2730_));
 sg13g2_nor2_1 _3674_ (.A(net460),
    .B(_2155_),
    .Y(_2732_));
 sg13g2_xnor2_1 _3675_ (.Y(_2733_),
    .A(net460),
    .B(_2154_));
 sg13g2_a21oi_1 _3676_ (.A1(_2694_),
    .A2(_2733_),
    .Y(_2735_),
    .B1(_2732_));
 sg13g2_xnor2_1 _3677_ (.Y(_2736_),
    .A(_2731_),
    .B(_2735_));
 sg13g2_xnor2_1 _3678_ (.Y(_2737_),
    .A(_2709_),
    .B(_2725_));
 sg13g2_nand2b_1 _3679_ (.Y(_2738_),
    .B(_2737_),
    .A_N(_2736_));
 sg13g2_o21ai_1 _3680_ (.B1(_2738_),
    .Y(_2739_),
    .A1(_2709_),
    .A2(_2726_));
 sg13g2_a21oi_1 _3681_ (.A1(_2703_),
    .A2(_2713_),
    .Y(_2740_),
    .B1(_2711_));
 sg13g2_nor2_1 _3682_ (.A(_2171_),
    .B(_2697_),
    .Y(_2741_));
 sg13g2_xor2_1 _3683_ (.B(_2697_),
    .A(_2171_),
    .X(_2742_));
 sg13g2_nor2b_1 _3684_ (.A(_2740_),
    .B_N(_2742_),
    .Y(_2743_));
 sg13g2_xnor2_1 _3685_ (.Y(_2744_),
    .A(_2740_),
    .B(_2742_));
 sg13g2_xor2_1 _3686_ (.B(_2744_),
    .A(_2727_),
    .X(_2746_));
 sg13g2_a21o_1 _3687_ (.A2(_2719_),
    .A1(_2632_),
    .B1(_2724_),
    .X(_2747_));
 sg13g2_nor3_1 _3688_ (.A(_2142_),
    .B(_2697_),
    .C(_2719_),
    .Y(_2748_));
 sg13g2_xnor2_1 _3689_ (.Y(_2749_),
    .A(_2697_),
    .B(_2721_));
 sg13g2_xnor2_1 _3690_ (.Y(_2750_),
    .A(_2171_),
    .B(_2716_));
 sg13g2_xnor2_1 _3691_ (.Y(_2751_),
    .A(_2749_),
    .B(_2750_));
 sg13g2_nor2b_1 _3692_ (.A(_2751_),
    .B_N(_2747_),
    .Y(_2752_));
 sg13g2_xnor2_1 _3693_ (.Y(_2753_),
    .A(_2747_),
    .B(_2751_));
 sg13g2_xor2_1 _3694_ (.B(_2753_),
    .A(_2746_),
    .X(_2754_));
 sg13g2_o21ai_1 _3695_ (.B1(_2729_),
    .Y(_2755_),
    .A1(_2731_),
    .A2(_2735_));
 sg13g2_xnor2_1 _3696_ (.Y(_0033_),
    .A(_2739_),
    .B(_2754_));
 sg13g2_nor2b_1 _3697_ (.A(_0033_),
    .B_N(_2755_),
    .Y(_0034_));
 sg13g2_a21oi_1 _3698_ (.A1(_2739_),
    .A2(_2754_),
    .Y(_0035_),
    .B1(_0034_));
 sg13g2_a21oi_1 _3699_ (.A1(_2727_),
    .A2(_2744_),
    .Y(_0036_),
    .B1(_2743_));
 sg13g2_a21o_1 _3700_ (.A2(_2753_),
    .A1(_2746_),
    .B1(_2752_),
    .X(_0037_));
 sg13g2_a21oi_1 _3701_ (.A1(_2677_),
    .A2(_2741_),
    .Y(_0038_),
    .B1(_2658_));
 sg13g2_a21o_1 _3702_ (.A2(_2750_),
    .A1(_2749_),
    .B1(_2748_),
    .X(_0039_));
 sg13g2_xnor2_1 _3703_ (.Y(_0040_),
    .A(net504),
    .B(_0039_));
 sg13g2_xnor2_1 _3704_ (.Y(_0041_),
    .A(_0038_),
    .B(_0040_));
 sg13g2_nand2_1 _3705_ (.Y(_0042_),
    .A(_0037_),
    .B(_0041_));
 sg13g2_xnor2_1 _3706_ (.Y(_0044_),
    .A(_0037_),
    .B(_0041_));
 sg13g2_xor2_1 _3707_ (.B(_0044_),
    .A(_0036_),
    .X(_0045_));
 sg13g2_nand2b_1 _3708_ (.Y(_0046_),
    .B(_0045_),
    .A_N(_0035_));
 sg13g2_xnor2_1 _3709_ (.Y(_0047_),
    .A(_0035_),
    .B(_0045_));
 sg13g2_xor2_1 _3710_ (.B(_2659_),
    .A(_2271_),
    .X(_0048_));
 sg13g2_nor2b_1 _3711_ (.A(_2266_),
    .B_N(_0048_),
    .Y(_0049_));
 sg13g2_nand2_1 _3712_ (.Y(_0050_),
    .A(net459),
    .B(net458));
 sg13g2_inv_1 _3713_ (.Y(_0051_),
    .A(_0050_));
 sg13g2_and3_2 _3714_ (.X(_0052_),
    .A(net459),
    .B(_2684_),
    .C(net458));
 sg13g2_nor2_1 _3715_ (.A(_2685_),
    .B(_0050_),
    .Y(_0053_));
 sg13g2_a22oi_1 _3716_ (.Y(_0055_),
    .B1(net458),
    .B2(_2666_),
    .A2(_2684_),
    .A1(net459));
 sg13g2_a21oi_1 _3717_ (.A1(_2666_),
    .A2(_0052_),
    .Y(_0056_),
    .B1(_0055_));
 sg13g2_xnor2_1 _3718_ (.Y(_0057_),
    .A(_2270_),
    .B(_0056_));
 sg13g2_xnor2_1 _3719_ (.Y(_0058_),
    .A(_2266_),
    .B(_0048_));
 sg13g2_a21oi_1 _3720_ (.A1(_0057_),
    .A2(_0058_),
    .Y(_0059_),
    .B1(_0049_));
 sg13g2_xnor2_1 _3721_ (.Y(_0060_),
    .A(_2687_),
    .B(_2688_));
 sg13g2_nor2_1 _3722_ (.A(_0059_),
    .B(_0060_),
    .Y(_0061_));
 sg13g2_xnor2_1 _3723_ (.Y(_0062_),
    .A(_2042_),
    .B(_2700_));
 sg13g2_xor2_1 _3724_ (.B(_0060_),
    .A(_0059_),
    .X(_0063_));
 sg13g2_a21oi_1 _3725_ (.A1(_0062_),
    .A2(_0063_),
    .Y(_0064_),
    .B1(_0061_));
 sg13g2_xnor2_1 _3726_ (.Y(_0066_),
    .A(_2692_),
    .B(_2708_));
 sg13g2_nor2_1 _3727_ (.A(_0064_),
    .B(_0066_),
    .Y(_0067_));
 sg13g2_xor2_1 _3728_ (.B(_0066_),
    .A(_0064_),
    .X(_0068_));
 sg13g2_a21o_1 _3729_ (.A2(_0056_),
    .A1(_2269_),
    .B1(_0053_),
    .X(_0069_));
 sg13g2_xnor2_1 _3730_ (.Y(_0070_),
    .A(_2693_),
    .B(_2733_));
 sg13g2_nand2_1 _3731_ (.Y(_0071_),
    .A(_0069_),
    .B(_0070_));
 sg13g2_xnor2_1 _3732_ (.Y(_0072_),
    .A(_0069_),
    .B(_0070_));
 sg13g2_xor2_1 _3733_ (.B(_0072_),
    .A(_2044_),
    .X(_0073_));
 sg13g2_a21oi_1 _3734_ (.A1(_0068_),
    .A2(_0073_),
    .Y(_0074_),
    .B1(_0067_));
 sg13g2_xnor2_1 _3735_ (.Y(_0075_),
    .A(_2736_),
    .B(_2737_));
 sg13g2_nor2b_1 _3736_ (.A(_0074_),
    .B_N(_0075_),
    .Y(_0077_));
 sg13g2_o21ai_1 _3737_ (.B1(_0071_),
    .Y(_0078_),
    .A1(_2044_),
    .A2(_0072_));
 sg13g2_xnor2_1 _3738_ (.Y(_0079_),
    .A(_0074_),
    .B(_0075_));
 sg13g2_a21oi_1 _3739_ (.A1(_0078_),
    .A2(_0079_),
    .Y(_0080_),
    .B1(_0077_));
 sg13g2_inv_1 _3740_ (.Y(_0081_),
    .A(_0080_));
 sg13g2_xor2_1 _3741_ (.B(_0033_),
    .A(_2755_),
    .X(_0082_));
 sg13g2_inv_1 _3742_ (.Y(_0083_),
    .A(_0082_));
 sg13g2_nand2_1 _3743_ (.Y(_0084_),
    .A(_0080_),
    .B(_0082_));
 sg13g2_nand2_1 _3744_ (.Y(_0085_),
    .A(_0081_),
    .B(_0083_));
 sg13g2_nand2_2 _3745_ (.Y(_0086_),
    .A(net649),
    .B(_2666_));
 sg13g2_nand4_1 _3746_ (.B(net648),
    .C(net498),
    .A(net600),
    .Y(_0088_),
    .D(net459));
 sg13g2_nand2_1 _3747_ (.Y(_0089_),
    .A(_2097_),
    .B(_0088_));
 sg13g2_a22oi_1 _3748_ (.Y(_0090_),
    .B1(net459),
    .B2(net648),
    .A2(net498),
    .A1(net600));
 sg13g2_a21o_1 _3749_ (.A2(_0088_),
    .A1(_2097_),
    .B1(_0090_),
    .X(_0091_));
 sg13g2_or2_1 _3750_ (.X(_0092_),
    .B(_0091_),
    .A(_0086_));
 sg13g2_xnor2_1 _3751_ (.Y(_0093_),
    .A(_0086_),
    .B(_0091_));
 sg13g2_nor2_1 _3752_ (.A(_2341_),
    .B(_0086_),
    .Y(_0094_));
 sg13g2_xor2_1 _3753_ (.B(_0086_),
    .A(_2341_),
    .X(_0095_));
 sg13g2_xnor2_1 _3754_ (.Y(_0096_),
    .A(_0051_),
    .B(_0095_));
 sg13g2_o21ai_1 _3755_ (.B1(_0092_),
    .Y(_0097_),
    .A1(_0093_),
    .A2(_0096_));
 sg13g2_xnor2_1 _3756_ (.Y(_0099_),
    .A(_0057_),
    .B(_0058_));
 sg13g2_nand2b_1 _3757_ (.Y(_0100_),
    .B(_0097_),
    .A_N(_0099_));
 sg13g2_xor2_1 _3758_ (.B(_0099_),
    .A(_0097_),
    .X(_0101_));
 sg13g2_a21oi_1 _3759_ (.A1(_0051_),
    .A2(_0095_),
    .Y(_0102_),
    .B1(_0094_));
 sg13g2_nor2b_1 _3760_ (.A(_0102_),
    .B_N(_0057_),
    .Y(_0103_));
 sg13g2_xnor2_1 _3761_ (.Y(_0104_),
    .A(_0057_),
    .B(_0102_));
 sg13g2_xnor2_1 _3762_ (.Y(_0105_),
    .A(_0052_),
    .B(_0104_));
 sg13g2_o21ai_1 _3763_ (.B1(_0100_),
    .Y(_0106_),
    .A1(_0101_),
    .A2(_0105_));
 sg13g2_xnor2_1 _3764_ (.Y(_0107_),
    .A(_0062_),
    .B(_0063_));
 sg13g2_nor2b_1 _3765_ (.A(_0107_),
    .B_N(_0106_),
    .Y(_0108_));
 sg13g2_nand2b_1 _3766_ (.Y(_0110_),
    .B(_0107_),
    .A_N(_0106_));
 sg13g2_nand2b_1 _3767_ (.Y(_0111_),
    .B(_0110_),
    .A_N(_0108_));
 sg13g2_a21oi_1 _3768_ (.A1(_0052_),
    .A2(_0104_),
    .Y(_0112_),
    .B1(_0103_));
 sg13g2_nor2b_1 _3769_ (.A(_0112_),
    .B_N(_2696_),
    .Y(_0113_));
 sg13g2_xnor2_1 _3770_ (.Y(_0114_),
    .A(_2696_),
    .B(_0112_));
 sg13g2_xor2_1 _3771_ (.B(_0114_),
    .A(_2660_),
    .X(_0115_));
 sg13g2_a21oi_1 _3772_ (.A1(_0110_),
    .A2(_0115_),
    .Y(_0116_),
    .B1(_0108_));
 sg13g2_xor2_1 _3773_ (.B(_0073_),
    .A(_0068_),
    .X(_0117_));
 sg13g2_nand2b_1 _3774_ (.Y(_0118_),
    .B(_0117_),
    .A_N(_0116_));
 sg13g2_a21o_1 _3775_ (.A2(_0114_),
    .A1(_2660_),
    .B1(_0113_),
    .X(_0119_));
 sg13g2_xnor2_1 _3776_ (.Y(_0121_),
    .A(_0116_),
    .B(_0117_));
 sg13g2_nand2_1 _3777_ (.Y(_0122_),
    .A(_0119_),
    .B(_0121_));
 sg13g2_xnor2_1 _3778_ (.Y(_0123_),
    .A(_0078_),
    .B(_0079_));
 sg13g2_nand3_1 _3779_ (.B(_0122_),
    .C(_0123_),
    .A(_0118_),
    .Y(_0124_));
 sg13g2_inv_1 _3780_ (.Y(_0125_),
    .A(_0124_));
 sg13g2_a21oi_1 _3781_ (.A1(_0118_),
    .A2(_0122_),
    .Y(_0126_),
    .B1(_0123_));
 sg13g2_xnor2_1 _3782_ (.Y(_0127_),
    .A(_0111_),
    .B(_0115_));
 sg13g2_and2_1 _3783_ (.A(net648),
    .B(_2684_),
    .X(_0128_));
 sg13g2_nand2_1 _3784_ (.Y(_0129_),
    .A(_1886_),
    .B(_0128_));
 sg13g2_nand3_1 _3785_ (.B(net501),
    .C(_0128_),
    .A(_1886_),
    .Y(_0130_));
 sg13g2_o21ai_1 _3786_ (.B1(_0130_),
    .Y(_0132_),
    .A1(_0089_),
    .A2(_0090_));
 sg13g2_xor2_1 _3787_ (.B(_0096_),
    .A(_0093_),
    .X(_0133_));
 sg13g2_nand2_1 _3788_ (.Y(_0134_),
    .A(_0132_),
    .B(_0133_));
 sg13g2_xnor2_1 _3789_ (.Y(_0135_),
    .A(_0132_),
    .B(_0133_));
 sg13g2_xor2_1 _3790_ (.B(_0050_),
    .A(_2684_),
    .X(_0136_));
 sg13g2_xor2_1 _3791_ (.B(_0136_),
    .A(_0088_),
    .X(_0137_));
 sg13g2_nand2b_1 _3792_ (.Y(_0138_),
    .B(_0137_),
    .A_N(_2698_));
 sg13g2_xor2_1 _3793_ (.B(_0137_),
    .A(_2698_),
    .X(_0139_));
 sg13g2_o21ai_1 _3794_ (.B1(_0134_),
    .Y(_0140_),
    .A1(_0135_),
    .A2(_0139_));
 sg13g2_xor2_1 _3795_ (.B(_0105_),
    .A(_0101_),
    .X(_0141_));
 sg13g2_nand2_1 _3796_ (.Y(_0143_),
    .A(_0140_),
    .B(_0141_));
 sg13g2_xnor2_1 _3797_ (.Y(_0144_),
    .A(_0140_),
    .B(_0141_));
 sg13g2_nand3_1 _3798_ (.B(net505),
    .C(net501),
    .A(net600),
    .Y(_0145_));
 sg13g2_o21ai_1 _3799_ (.B1(_0138_),
    .Y(_0146_),
    .A1(_0088_),
    .A2(_0136_));
 sg13g2_xor2_1 _3800_ (.B(_0146_),
    .A(_0048_),
    .X(_0147_));
 sg13g2_nor2b_1 _3801_ (.A(_0145_),
    .B_N(_0147_),
    .Y(_0148_));
 sg13g2_xor2_1 _3802_ (.B(_0147_),
    .A(_0145_),
    .X(_0149_));
 sg13g2_o21ai_1 _3803_ (.B1(_0143_),
    .Y(_0150_),
    .A1(_0144_),
    .A2(_0149_));
 sg13g2_nand2_1 _3804_ (.Y(_0151_),
    .A(_0127_),
    .B(_0150_));
 sg13g2_a21oi_1 _3805_ (.A1(_0048_),
    .A2(_0146_),
    .Y(_0152_),
    .B1(_0148_));
 sg13g2_xnor2_1 _3806_ (.Y(_0154_),
    .A(_0127_),
    .B(_0150_));
 sg13g2_o21ai_1 _3807_ (.B1(_0151_),
    .Y(_0155_),
    .A1(_0152_),
    .A2(_0154_));
 sg13g2_xor2_1 _3808_ (.B(_0121_),
    .A(_0119_),
    .X(_0156_));
 sg13g2_nand2_1 _3809_ (.Y(_0157_),
    .A(_0155_),
    .B(_0156_));
 sg13g2_a22oi_1 _3810_ (.Y(_0158_),
    .B1(_0129_),
    .B2(_2097_),
    .A2(_0128_),
    .A1(net501));
 sg13g2_nand4_1 _3811_ (.B(net648),
    .C(_1853_),
    .A(net600),
    .Y(_0159_),
    .D(net458));
 sg13g2_xnor2_1 _3812_ (.Y(_0160_),
    .A(_1897_),
    .B(_0128_));
 sg13g2_nor2b_1 _3813_ (.A(_0159_),
    .B_N(_0160_),
    .Y(_0161_));
 sg13g2_xnor2_1 _3814_ (.Y(_0162_),
    .A(_0159_),
    .B(_0160_));
 sg13g2_a21oi_1 _3815_ (.A1(_2422_),
    .A2(_0162_),
    .Y(_0163_),
    .B1(_0161_));
 sg13g2_nand2b_1 _3816_ (.Y(_0165_),
    .B(_0158_),
    .A_N(_0163_));
 sg13g2_nand2_1 _3817_ (.Y(_0166_),
    .A(_2695_),
    .B(_0128_));
 sg13g2_xor2_1 _3818_ (.B(_0163_),
    .A(_0158_),
    .X(_0167_));
 sg13g2_o21ai_1 _3819_ (.B1(_0165_),
    .Y(_0168_),
    .A1(_0166_),
    .A2(_0167_));
 sg13g2_xor2_1 _3820_ (.B(_0139_),
    .A(_0135_),
    .X(_0169_));
 sg13g2_xnor2_1 _3821_ (.Y(_0170_),
    .A(_2039_),
    .B(_2341_));
 sg13g2_inv_1 _3822_ (.Y(_0171_),
    .A(_0170_));
 sg13g2_xnor2_1 _3823_ (.Y(_0172_),
    .A(_0168_),
    .B(_0169_));
 sg13g2_nor2_1 _3824_ (.A(_0170_),
    .B(_0172_),
    .Y(_0173_));
 sg13g2_nand2_1 _3825_ (.Y(_0174_),
    .A(_0170_),
    .B(_0172_));
 sg13g2_nand3_1 _3826_ (.B(_2422_),
    .C(net458),
    .A(net648),
    .Y(_0176_));
 sg13g2_a21oi_1 _3827_ (.A1(net653),
    .A2(_2695_),
    .Y(_0177_),
    .B1(_1875_));
 sg13g2_xor2_1 _3828_ (.B(_0162_),
    .A(_2422_),
    .X(_0178_));
 sg13g2_nand2_1 _3829_ (.Y(_0179_),
    .A(_0177_),
    .B(_0178_));
 sg13g2_xnor2_1 _3830_ (.Y(_0180_),
    .A(_0177_),
    .B(_0178_));
 sg13g2_o21ai_1 _3831_ (.B1(_2647_),
    .Y(_0181_),
    .A1(net648),
    .A2(_2668_));
 sg13g2_a21oi_1 _3832_ (.A1(net648),
    .A2(net458),
    .Y(_0182_),
    .B1(_2422_));
 sg13g2_xnor2_1 _3833_ (.Y(_0183_),
    .A(_0180_),
    .B(_0181_));
 sg13g2_a21oi_1 _3834_ (.A1(_0176_),
    .A2(_0183_),
    .Y(_0184_),
    .B1(_0182_));
 sg13g2_xor2_1 _3835_ (.B(_0167_),
    .A(_0166_),
    .X(_0185_));
 sg13g2_o21ai_1 _3836_ (.B1(_0179_),
    .Y(_0187_),
    .A1(_0180_),
    .A2(_0181_));
 sg13g2_a21oi_1 _3837_ (.A1(_2096_),
    .A2(_0187_),
    .Y(_0188_),
    .B1(_0185_));
 sg13g2_nor2b_1 _3838_ (.A(_0184_),
    .B_N(_0188_),
    .Y(_0189_));
 sg13g2_a221oi_1 _3839_ (.B2(_0185_),
    .C1(_0187_),
    .B1(_0184_),
    .A1(_1886_),
    .Y(_0190_),
    .A2(net501));
 sg13g2_nor2_1 _3840_ (.A(_0189_),
    .B(_0190_),
    .Y(_0191_));
 sg13g2_nand4_1 _3841_ (.B(_0169_),
    .C(_0171_),
    .A(_0168_),
    .Y(_0192_),
    .D(_0191_));
 sg13g2_xnor2_1 _3842_ (.Y(_0193_),
    .A(_0144_),
    .B(_0149_));
 sg13g2_a221oi_1 _3843_ (.B2(_0191_),
    .C1(_0173_),
    .B1(_0174_),
    .A1(_0168_),
    .Y(_0194_),
    .A2(_0169_));
 sg13g2_a221oi_1 _3844_ (.B2(_0193_),
    .C1(_0194_),
    .B1(_0192_),
    .A1(_0152_),
    .Y(_0195_),
    .A2(_0154_));
 sg13g2_o21ai_1 _3845_ (.B1(_0195_),
    .Y(_0196_),
    .A1(_0152_),
    .A2(_0154_));
 sg13g2_xnor2_1 _3846_ (.Y(_0198_),
    .A(_0155_),
    .B(_0156_));
 sg13g2_o21ai_1 _3847_ (.B1(_0157_),
    .Y(_0199_),
    .A1(_0196_),
    .A2(_0198_));
 sg13g2_nor2_1 _3848_ (.A(_0125_),
    .B(_0126_),
    .Y(_0200_));
 sg13g2_a221oi_1 _3849_ (.B2(_0199_),
    .C1(_0126_),
    .B1(_0124_),
    .A1(_0081_),
    .Y(_0201_),
    .A2(_0083_));
 sg13g2_a21oi_2 _3850_ (.B1(_0201_),
    .Y(_0202_),
    .A2(_0082_),
    .A1(_0080_));
 sg13g2_nand2_1 _3851_ (.Y(_0203_),
    .A(_0047_),
    .B(_0202_));
 sg13g2_o21ai_1 _3852_ (.B1(_0042_),
    .Y(_0204_),
    .A1(_0036_),
    .A2(_0044_));
 sg13g2_a21oi_1 _3853_ (.A1(net504),
    .A2(_0038_),
    .Y(_0205_),
    .B1(_0039_));
 sg13g2_nor2_1 _3854_ (.A(_2741_),
    .B(_0205_),
    .Y(_0206_));
 sg13g2_xnor2_1 _3855_ (.Y(_0207_),
    .A(_0204_),
    .B(_0206_));
 sg13g2_a21o_1 _3856_ (.A2(_0203_),
    .A1(_0046_),
    .B1(_0207_),
    .X(_0209_));
 sg13g2_nand3_1 _3857_ (.B(_0203_),
    .C(_0207_),
    .A(_0046_),
    .Y(_0210_));
 sg13g2_a221oi_1 _3858_ (.B2(_0200_),
    .C1(_0126_),
    .B1(_0199_),
    .A1(_0084_),
    .Y(_0211_),
    .A2(_0085_));
 sg13g2_nor2_1 _3859_ (.A(_0199_),
    .B(_0200_),
    .Y(_0212_));
 sg13g2_xnor2_1 _3860_ (.Y(_0213_),
    .A(_0196_),
    .B(_0198_));
 sg13g2_nor3_2 _3861_ (.A(_0211_),
    .B(_0212_),
    .C(_0213_),
    .Y(_0214_));
 sg13g2_a21oi_1 _3862_ (.A1(net600),
    .A2(net536),
    .Y(_0215_),
    .B1(net650));
 sg13g2_o21ai_1 _3863_ (.B1(_0215_),
    .Y(_0216_),
    .A1(net600),
    .A2(net536));
 sg13g2_a21o_1 _3864_ (.A2(_1853_),
    .A1(net646),
    .B1(_0216_),
    .X(_0217_));
 sg13g2_o21ai_1 _3865_ (.B1(_0217_),
    .Y(_0218_),
    .A1(net646),
    .A2(_1853_));
 sg13g2_o21ai_1 _3866_ (.B1(_0218_),
    .Y(_0220_),
    .A1(net641),
    .A2(_2420_));
 sg13g2_nor2_2 _3867_ (.A(_0736_),
    .B(_2667_),
    .Y(_0221_));
 sg13g2_inv_1 _3868_ (.Y(_0222_),
    .A(_0221_));
 sg13g2_a22oi_1 _3869_ (.Y(_0223_),
    .B1(_0221_),
    .B2(_2329_),
    .A2(_2420_),
    .A1(net641));
 sg13g2_a21oi_2 _3870_ (.B1(_1120_),
    .Y(_0224_),
    .A2(_1109_),
    .A1(net589));
 sg13g2_nand2b_2 _3871_ (.Y(_0225_),
    .B(_2025_),
    .A_N(_1120_));
 sg13g2_nor2_2 _3872_ (.A(net640),
    .B(_0945_),
    .Y(_0226_));
 sg13g2_xnor2_1 _3873_ (.Y(_0227_),
    .A(net633),
    .B(_0736_));
 sg13g2_a22oi_1 _3874_ (.Y(_0228_),
    .B1(_0223_),
    .B2(_0220_),
    .A2(_0222_),
    .A1(net497));
 sg13g2_o21ai_1 _3875_ (.B1(_0228_),
    .Y(_0229_),
    .A1(net476),
    .A2(_0227_));
 sg13g2_xnor2_1 _3876_ (.Y(_0231_),
    .A(net626),
    .B(_0226_));
 sg13g2_a22oi_1 _3877_ (.Y(_0232_),
    .B1(_0231_),
    .B2(net584),
    .A2(_0227_),
    .A1(net476));
 sg13g2_a21oi_2 _3878_ (.B1(net556),
    .Y(_0233_),
    .A2(_0912_),
    .A1(_0736_));
 sg13g2_nor2_2 _3879_ (.A(net627),
    .B(net621),
    .Y(_0234_));
 sg13g2_inv_2 _3880_ (.Y(_0235_),
    .A(_0234_));
 sg13g2_a21oi_1 _3881_ (.A1(_0226_),
    .A2(_0234_),
    .Y(_0236_),
    .B1(_0233_));
 sg13g2_nor2_1 _3882_ (.A(net567),
    .B(net578),
    .Y(_0237_));
 sg13g2_nor2_2 _3883_ (.A(_0516_),
    .B(_2572_),
    .Y(_0238_));
 sg13g2_a21oi_2 _3884_ (.B1(_0237_),
    .Y(_0239_),
    .A2(_0238_),
    .A1(net567));
 sg13g2_a21o_2 _3885_ (.A2(_0238_),
    .A1(net567),
    .B1(_0237_),
    .X(_0240_));
 sg13g2_nor2_1 _3886_ (.A(net584),
    .B(_0231_),
    .Y(_0242_));
 sg13g2_a221oi_1 _3887_ (.B2(_0240_),
    .C1(_0242_),
    .B1(_0236_),
    .A1(_0229_),
    .Y(_0243_),
    .A2(_0232_));
 sg13g2_and2_1 _3888_ (.A(_0549_),
    .B(_2605_),
    .X(_0244_));
 sg13g2_a21oi_2 _3889_ (.B1(net541),
    .Y(_0245_),
    .A2(_0244_),
    .A1(net570));
 sg13g2_a21o_2 _3890_ (.A2(_0244_),
    .A1(net570),
    .B1(net541),
    .X(_0246_));
 sg13g2_o21ai_1 _3891_ (.B1(_0245_),
    .Y(_0247_),
    .A1(net554),
    .A2(_0233_));
 sg13g2_a21o_1 _3892_ (.A2(_0233_),
    .A1(net554),
    .B1(_0247_),
    .X(_0248_));
 sg13g2_o21ai_1 _3893_ (.B1(_0248_),
    .Y(_0249_),
    .A1(_0236_),
    .A2(_0240_));
 sg13g2_nor2_2 _3894_ (.A(net616),
    .B(_0246_),
    .Y(_0250_));
 sg13g2_inv_1 _3895_ (.Y(_0251_),
    .A(_0250_));
 sg13g2_o21ai_1 _3896_ (.B1(_1755_),
    .Y(_0253_),
    .A1(net554),
    .A2(_0245_));
 sg13g2_a21oi_1 _3897_ (.A1(_0233_),
    .A2(_0251_),
    .Y(_0254_),
    .B1(_0253_));
 sg13g2_o21ai_1 _3898_ (.B1(_0254_),
    .Y(_0255_),
    .A1(_0243_),
    .A2(_0249_));
 sg13g2_nand3_1 _3899_ (.B(_2329_),
    .C(net476),
    .A(net585),
    .Y(_0256_));
 sg13g2_o21ai_1 _3900_ (.B1(_0240_),
    .Y(_0257_),
    .A1(net580),
    .A2(_0256_));
 sg13g2_nand2_1 _3901_ (.Y(_0258_),
    .A(_0648_),
    .B(_1755_));
 sg13g2_o21ai_1 _3902_ (.B1(_0257_),
    .Y(_0259_),
    .A1(_0923_),
    .A2(_0258_));
 sg13g2_nor4_2 _3903_ (.A(_0214_),
    .B(_0246_),
    .C(_0255_),
    .Y(_0260_),
    .D(_0259_));
 sg13g2_xnor2_1 _3904_ (.Y(_0261_),
    .A(_0047_),
    .B(_0202_));
 sg13g2_nand4_1 _3905_ (.B(_0210_),
    .C(_0260_),
    .A(_0209_),
    .Y(_0262_),
    .D(_0261_));
 sg13g2_nor2_2 _3906_ (.A(net550),
    .B(_0428_),
    .Y(_0264_));
 sg13g2_nand2b_1 _3907_ (.Y(_0265_),
    .B(_0417_),
    .A_N(net550));
 sg13g2_and2_1 _3908_ (.A(_0263_),
    .B(_0439_),
    .X(_0266_));
 sg13g2_nand2_2 _3909_ (.Y(_0267_),
    .A(_0263_),
    .B(_0439_));
 sg13g2_nor2_1 _3910_ (.A(net473),
    .B(_0267_),
    .Y(_0268_));
 sg13g2_nand2_1 _3911_ (.Y(_0269_),
    .A(_0264_),
    .B(_0266_));
 sg13g2_nor2_2 _3912_ (.A(net585),
    .B(net476),
    .Y(_0270_));
 sg13g2_nand2_1 _3913_ (.Y(_0271_),
    .A(net497),
    .B(_0270_));
 sg13g2_nand2_1 _3914_ (.Y(_0272_),
    .A(net497),
    .B(_2421_));
 sg13g2_nor2_1 _3915_ (.A(_2420_),
    .B(_0271_),
    .Y(_0273_));
 sg13g2_o21ai_1 _3916_ (.B1(net475),
    .Y(_0275_),
    .A1(_2420_),
    .A2(_0271_));
 sg13g2_a21o_1 _3917_ (.A2(_0275_),
    .A1(_0251_),
    .B1(_0253_),
    .X(_0276_));
 sg13g2_nand2_1 _3918_ (.Y(_0277_),
    .A(net637),
    .B(_2448_));
 sg13g2_o21ai_1 _3919_ (.B1(_0218_),
    .Y(_0278_),
    .A1(_2690_),
    .A2(_2421_));
 sg13g2_o21ai_1 _3920_ (.B1(_0278_),
    .Y(_0279_),
    .A1(net641),
    .A2(_2420_));
 sg13g2_xnor2_1 _3921_ (.Y(_0280_),
    .A(_0225_),
    .B(_0272_));
 sg13g2_nand2_1 _3922_ (.Y(_0281_),
    .A(net558),
    .B(_2449_));
 sg13g2_o21ai_1 _3923_ (.B1(_0281_),
    .Y(_0282_),
    .A1(net633),
    .A2(_0280_));
 sg13g2_a21oi_1 _3924_ (.A1(_0277_),
    .A2(_0279_),
    .Y(_0283_),
    .B1(_0282_));
 sg13g2_o21ai_1 _3925_ (.B1(net585),
    .Y(_0284_),
    .A1(net476),
    .A2(_0272_));
 sg13g2_nor2b_1 _3926_ (.A(_0273_),
    .B_N(_0284_),
    .Y(_0286_));
 sg13g2_a221oi_1 _3927_ (.B2(net626),
    .C1(_0283_),
    .B1(_0286_),
    .A1(net633),
    .Y(_0287_),
    .A2(_0280_));
 sg13g2_nand2_2 _3928_ (.Y(_0288_),
    .A(_0240_),
    .B(_0270_));
 sg13g2_nor2_1 _3929_ (.A(_2329_),
    .B(_0288_),
    .Y(_0289_));
 sg13g2_o21ai_1 _3930_ (.B1(_0275_),
    .Y(_0290_),
    .A1(_0272_),
    .A2(_0288_));
 sg13g2_or2_1 _3931_ (.X(_0291_),
    .B(_0286_),
    .A(net626));
 sg13g2_o21ai_1 _3932_ (.B1(_0291_),
    .Y(_0292_),
    .A1(net621),
    .A2(_0290_));
 sg13g2_nand2b_1 _3933_ (.Y(_0293_),
    .B(net551),
    .A_N(_0275_));
 sg13g2_nor2_1 _3934_ (.A(net614),
    .B(_0245_),
    .Y(_0294_));
 sg13g2_nor3_1 _3935_ (.A(_0250_),
    .B(_0275_),
    .C(_0294_),
    .Y(_0295_));
 sg13g2_a22oi_1 _3936_ (.Y(_0297_),
    .B1(_0293_),
    .B2(_0253_),
    .A2(_0290_),
    .A1(net621));
 sg13g2_o21ai_1 _3937_ (.B1(_0297_),
    .Y(_0298_),
    .A1(_0287_),
    .A2(_0292_));
 sg13g2_o21ai_1 _3938_ (.B1(_0276_),
    .Y(_0299_),
    .A1(_0295_),
    .A2(_0298_));
 sg13g2_inv_1 _3939_ (.Y(_0300_),
    .A(_0299_));
 sg13g2_xnor2_1 _3940_ (.Y(_0301_),
    .A(net634),
    .B(_0224_));
 sg13g2_inv_1 _3941_ (.Y(_0302_),
    .A(_0301_));
 sg13g2_nor2_1 _3942_ (.A(net641),
    .B(_2421_),
    .Y(_0303_));
 sg13g2_nand2_1 _3943_ (.Y(_0304_),
    .A(net641),
    .B(_2421_));
 sg13g2_o21ai_1 _3944_ (.B1(_0304_),
    .Y(_0305_),
    .A1(_0218_),
    .A2(_0303_));
 sg13g2_a21oi_1 _3945_ (.A1(net637),
    .A2(net497),
    .Y(_0306_),
    .B1(_0305_));
 sg13g2_a21oi_1 _3946_ (.A1(net558),
    .A2(_2329_),
    .Y(_0308_),
    .B1(_0306_));
 sg13g2_nor2b_1 _3947_ (.A(net585),
    .B_N(net628),
    .Y(_0309_));
 sg13g2_nor2_1 _3948_ (.A(_2580_),
    .B(net628),
    .Y(_0310_));
 sg13g2_nor3_1 _3949_ (.A(_0302_),
    .B(_0309_),
    .C(_0310_),
    .Y(_0311_));
 sg13g2_xnor2_1 _3950_ (.Y(_0312_),
    .A(_2580_),
    .B(net476));
 sg13g2_a221oi_1 _3951_ (.B2(net626),
    .C1(_0311_),
    .B1(_0312_),
    .A1(_0302_),
    .Y(_0313_),
    .A2(_0308_));
 sg13g2_or2_1 _3952_ (.X(_0314_),
    .B(_0312_),
    .A(net628));
 sg13g2_xnor2_1 _3953_ (.Y(_0315_),
    .A(_0239_),
    .B(_0270_));
 sg13g2_o21ai_1 _3954_ (.B1(_0314_),
    .Y(_0316_),
    .A1(net622),
    .A2(_0315_));
 sg13g2_nor2_1 _3955_ (.A(_0245_),
    .B(_0288_),
    .Y(_0317_));
 sg13g2_xnor2_1 _3956_ (.Y(_0319_),
    .A(_0246_),
    .B(_0288_));
 sg13g2_a22oi_1 _3957_ (.Y(_0320_),
    .B1(_0319_),
    .B2(net616),
    .A2(_0315_),
    .A1(net622));
 sg13g2_o21ai_1 _3958_ (.B1(_0320_),
    .Y(_0321_),
    .A1(_0313_),
    .A2(_0316_));
 sg13g2_nor2_1 _3959_ (.A(net616),
    .B(_0319_),
    .Y(_0322_));
 sg13g2_nor2_1 _3960_ (.A(net611),
    .B(_0317_),
    .Y(_0323_));
 sg13g2_nor2_1 _3961_ (.A(_0322_),
    .B(_0323_),
    .Y(_0324_));
 sg13g2_a221oi_1 _3962_ (.B2(_0324_),
    .C1(net606),
    .B1(_0321_),
    .A1(net611),
    .Y(_0325_),
    .A2(_0317_));
 sg13g2_o21ai_1 _3963_ (.B1(_0300_),
    .Y(_0326_),
    .A1(net538),
    .A2(_0325_));
 sg13g2_nand3_1 _3964_ (.B(_0268_),
    .C(_0326_),
    .A(_0262_),
    .Y(_0327_));
 sg13g2_nand3_1 _3965_ (.B(_0296_),
    .C(_2565_),
    .A(_0153_),
    .Y(_0328_));
 sg13g2_inv_1 _3966_ (.Y(_0330_),
    .A(_0328_));
 sg13g2_nor2_2 _3967_ (.A(net618),
    .B(net553),
    .Y(_0331_));
 sg13g2_nor2_1 _3968_ (.A(_2620_),
    .B(_0331_),
    .Y(_0332_));
 sg13g2_nor2b_1 _3969_ (.A(net621),
    .B_N(net627),
    .Y(_0333_));
 sg13g2_xor2_1 _3970_ (.B(net622),
    .A(net629),
    .X(_0334_));
 sg13g2_nor2_2 _3971_ (.A(_2643_),
    .B(_2678_),
    .Y(_0335_));
 sg13g2_a21oi_2 _3972_ (.B1(_1427_),
    .Y(_0336_),
    .A2(_0335_),
    .A1(_0945_));
 sg13g2_a21oi_1 _3973_ (.A1(_2557_),
    .A2(_0336_),
    .Y(_0337_),
    .B1(_0912_));
 sg13g2_a21oi_1 _3974_ (.A1(_0334_),
    .A2(_0337_),
    .Y(_0338_),
    .B1(_2637_));
 sg13g2_a21oi_2 _3975_ (.B1(_0648_),
    .Y(_0339_),
    .A2(_0338_),
    .A1(_2553_));
 sg13g2_nand2b_1 _3976_ (.Y(_0341_),
    .B(_0339_),
    .A_N(_0332_));
 sg13g2_xor2_1 _3977_ (.B(_0339_),
    .A(_0332_),
    .X(_0342_));
 sg13g2_nor2_1 _3978_ (.A(net581),
    .B(_0342_),
    .Y(_0343_));
 sg13g2_xor2_1 _3979_ (.B(net607),
    .A(net612),
    .X(_0344_));
 sg13g2_nand2_1 _3980_ (.Y(_0345_),
    .A(_2594_),
    .B(_0341_));
 sg13g2_xnor2_1 _3981_ (.Y(_0346_),
    .A(_0344_),
    .B(_0345_));
 sg13g2_nand2_1 _3982_ (.Y(_0347_),
    .A(net575),
    .B(_0346_));
 sg13g2_xnor2_1 _3983_ (.Y(_0348_),
    .A(net575),
    .B(_0346_));
 sg13g2_nand2_1 _3984_ (.Y(_0349_),
    .A(_0343_),
    .B(_0348_));
 sg13g2_xor2_1 _3985_ (.B(_0338_),
    .A(_1744_),
    .X(_0350_));
 sg13g2_nor2_1 _3986_ (.A(net586),
    .B(_0350_),
    .Y(_0352_));
 sg13g2_xor2_1 _3987_ (.B(_0342_),
    .A(net581),
    .X(_0353_));
 sg13g2_xnor2_1 _3988_ (.Y(_0354_),
    .A(_0352_),
    .B(_0353_));
 sg13g2_xnor2_1 _3989_ (.Y(_0355_),
    .A(_0334_),
    .B(_0337_));
 sg13g2_nand2_1 _3990_ (.Y(_0356_),
    .A(net591),
    .B(_0355_));
 sg13g2_xnor2_1 _3991_ (.Y(_0357_),
    .A(_2580_),
    .B(_0350_));
 sg13g2_nor2_1 _3992_ (.A(_0356_),
    .B(_0357_),
    .Y(_0358_));
 sg13g2_nor2_1 _3993_ (.A(net557),
    .B(net626),
    .Y(_0359_));
 sg13g2_xnor2_1 _3994_ (.Y(_0360_),
    .A(net635),
    .B(net631));
 sg13g2_xnor2_1 _3995_ (.Y(_0361_),
    .A(_0336_),
    .B(_0360_));
 sg13g2_nor2_2 _3996_ (.A(net592),
    .B(_0361_),
    .Y(_0363_));
 sg13g2_inv_1 _3997_ (.Y(_0364_),
    .A(_0363_));
 sg13g2_xnor2_1 _3998_ (.Y(_0365_),
    .A(_2591_),
    .B(_0355_));
 sg13g2_xnor2_1 _3999_ (.Y(_0366_),
    .A(_1438_),
    .B(_0335_));
 sg13g2_nand2_1 _4000_ (.Y(_0367_),
    .A(net597),
    .B(_0366_));
 sg13g2_xnor2_1 _4001_ (.Y(_0368_),
    .A(net561),
    .B(_0361_));
 sg13g2_o21ai_1 _4002_ (.B1(net645),
    .Y(_0369_),
    .A1(net650),
    .A2(net640));
 sg13g2_xor2_1 _4003_ (.B(_0369_),
    .A(_0221_),
    .X(_0370_));
 sg13g2_xnor2_1 _4004_ (.Y(_0371_),
    .A(_2613_),
    .B(_0366_));
 sg13g2_a21oi_1 _4005_ (.A1(net598),
    .A2(_0370_),
    .Y(_0372_),
    .B1(_0371_));
 sg13g2_o21ai_1 _4006_ (.B1(_2647_),
    .Y(_0374_),
    .A1(net649),
    .A2(_2683_));
 sg13g2_nor2_1 _4007_ (.A(_2635_),
    .B(_0374_),
    .Y(_0375_));
 sg13g2_xnor2_1 _4008_ (.Y(_0376_),
    .A(_2624_),
    .B(_0370_));
 sg13g2_nor2_1 _4009_ (.A(_0375_),
    .B(_0376_),
    .Y(_0377_));
 sg13g2_nand3_1 _4010_ (.B(_0370_),
    .C(_0371_),
    .A(net598),
    .Y(_0378_));
 sg13g2_nor2b_1 _4011_ (.A(_0372_),
    .B_N(_0378_),
    .Y(_0379_));
 sg13g2_a21o_1 _4012_ (.A2(_0379_),
    .A1(_0377_),
    .B1(_0372_),
    .X(_0380_));
 sg13g2_xnor2_1 _4013_ (.Y(_0381_),
    .A(_0367_),
    .B(_0368_));
 sg13g2_nor2b_1 _4014_ (.A(_0381_),
    .B_N(_0380_),
    .Y(_0382_));
 sg13g2_a21o_2 _4015_ (.A2(_0368_),
    .A1(_0367_),
    .B1(_0382_),
    .X(_0383_));
 sg13g2_xnor2_1 _4016_ (.Y(_0385_),
    .A(_0363_),
    .B(_0365_));
 sg13g2_nand2_1 _4017_ (.Y(_0386_),
    .A(_0383_),
    .B(_0385_));
 sg13g2_o21ai_1 _4018_ (.B1(_0386_),
    .Y(_0387_),
    .A1(_0364_),
    .A2(_0365_));
 sg13g2_a21oi_1 _4019_ (.A1(_0356_),
    .A2(_0357_),
    .Y(_0388_),
    .B1(_0387_));
 sg13g2_nor2_1 _4020_ (.A(_0358_),
    .B(_0388_),
    .Y(_0389_));
 sg13g2_nor3_1 _4021_ (.A(_0354_),
    .B(_0358_),
    .C(_0388_),
    .Y(_0390_));
 sg13g2_a21o_1 _4022_ (.A2(_0353_),
    .A1(_0352_),
    .B1(_0390_),
    .X(_0391_));
 sg13g2_xor2_1 _4023_ (.B(_0348_),
    .A(_0343_),
    .X(_0392_));
 sg13g2_nand2_1 _4024_ (.Y(_0393_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_nand2_1 _4025_ (.Y(_0394_),
    .A(_0349_),
    .B(_0393_));
 sg13g2_nor3_1 _4026_ (.A(net618),
    .B(net607),
    .C(_0339_),
    .Y(_0396_));
 sg13g2_nor2_1 _4027_ (.A(_1755_),
    .B(_0396_),
    .Y(_0397_));
 sg13g2_inv_1 _4028_ (.Y(_0398_),
    .A(_0397_));
 sg13g2_o21ai_1 _4029_ (.B1(_0626_),
    .Y(_0399_),
    .A1(net612),
    .A2(_0339_));
 sg13g2_nand2_1 _4030_ (.Y(_0400_),
    .A(_0397_),
    .B(_0399_));
 sg13g2_xnor2_1 _4031_ (.Y(_0401_),
    .A(net565),
    .B(_0400_));
 sg13g2_xnor2_1 _4032_ (.Y(_0402_),
    .A(_0347_),
    .B(_0401_));
 sg13g2_a21oi_1 _4033_ (.A1(_0349_),
    .A2(_0393_),
    .Y(_0403_),
    .B1(_0402_));
 sg13g2_xor2_1 _4034_ (.B(_0402_),
    .A(_0394_),
    .X(_0404_));
 sg13g2_o21ai_1 _4035_ (.B1(_0399_),
    .Y(_0405_),
    .A1(net571),
    .A2(_0398_));
 sg13g2_a21o_1 _4036_ (.A2(_0401_),
    .A1(_0347_),
    .B1(_0403_),
    .X(_0407_));
 sg13g2_xor2_1 _4037_ (.B(_0407_),
    .A(_0405_),
    .X(_0408_));
 sg13g2_and2_1 _4038_ (.A(_0404_),
    .B(_0408_),
    .X(_0409_));
 sg13g2_xnor2_1 _4039_ (.Y(_0410_),
    .A(_0377_),
    .B(_0379_));
 sg13g2_xor2_1 _4040_ (.B(_0381_),
    .A(_0380_),
    .X(_0411_));
 sg13g2_nand2_1 _4041_ (.Y(_0412_),
    .A(_0410_),
    .B(_0411_));
 sg13g2_xnor2_1 _4042_ (.Y(_0413_),
    .A(_0356_),
    .B(_0357_));
 sg13g2_xnor2_1 _4043_ (.Y(_0414_),
    .A(_0387_),
    .B(_0413_));
 sg13g2_or2_1 _4044_ (.X(_0415_),
    .B(_0385_),
    .A(_0383_));
 sg13g2_and3_2 _4045_ (.X(_0416_),
    .A(_0386_),
    .B(_0414_),
    .C(_0415_));
 sg13g2_xnor2_1 _4046_ (.Y(_0418_),
    .A(_0354_),
    .B(_0389_));
 sg13g2_a21oi_1 _4047_ (.A1(_0412_),
    .A2(_0416_),
    .Y(_0419_),
    .B1(_0418_));
 sg13g2_xnor2_1 _4048_ (.Y(_0420_),
    .A(_0391_),
    .B(_0392_));
 sg13g2_o21ai_1 _4049_ (.B1(_0409_),
    .Y(_0421_),
    .A1(_0419_),
    .A2(_0420_));
 sg13g2_nand2_1 _4050_ (.Y(_0422_),
    .A(_0330_),
    .B(_0421_));
 sg13g2_a21oi_1 _4051_ (.A1(net601),
    .A2(_1021_),
    .Y(_0423_),
    .B1(net598));
 sg13g2_nor2_1 _4052_ (.A(_0374_),
    .B(_0423_),
    .Y(_0424_));
 sg13g2_nor2_2 _4053_ (.A(_2624_),
    .B(_2635_),
    .Y(_0425_));
 sg13g2_nand2_1 _4054_ (.Y(_0426_),
    .A(net598),
    .B(net601));
 sg13g2_a221oi_1 _4055_ (.B2(_1021_),
    .C1(_0424_),
    .B1(_0425_),
    .A1(net595),
    .Y(_0427_),
    .A2(_0370_));
 sg13g2_nand2b_1 _4056_ (.Y(_0429_),
    .B(net561),
    .A_N(_0366_));
 sg13g2_o21ai_1 _4057_ (.B1(_0429_),
    .Y(_0430_),
    .A1(net595),
    .A2(_0370_));
 sg13g2_a22oi_1 _4058_ (.Y(_0431_),
    .B1(_0366_),
    .B2(net592),
    .A2(_0361_),
    .A1(net587));
 sg13g2_o21ai_1 _4059_ (.B1(_0431_),
    .Y(_0432_),
    .A1(_0427_),
    .A2(_0430_));
 sg13g2_nor2_1 _4060_ (.A(net585),
    .B(_0355_),
    .Y(_0433_));
 sg13g2_o21ai_1 _4061_ (.B1(_0432_),
    .Y(_0434_),
    .A1(net587),
    .A2(_0361_));
 sg13g2_a22oi_1 _4062_ (.Y(_0435_),
    .B1(_0355_),
    .B2(net586),
    .A2(_0350_),
    .A1(net580));
 sg13g2_o21ai_1 _4063_ (.B1(_0435_),
    .Y(_0436_),
    .A1(_0433_),
    .A2(_0434_));
 sg13g2_nor2_1 _4064_ (.A(net575),
    .B(_0342_),
    .Y(_0437_));
 sg13g2_o21ai_1 _4065_ (.B1(_0436_),
    .Y(_0438_),
    .A1(net581),
    .A2(_0350_));
 sg13g2_a22oi_1 _4066_ (.Y(_0440_),
    .B1(_0346_),
    .B2(net571),
    .A2(_0342_),
    .A1(net575));
 sg13g2_o21ai_1 _4067_ (.B1(_0440_),
    .Y(_0441_),
    .A1(_0437_),
    .A2(_0438_));
 sg13g2_o21ai_1 _4068_ (.B1(_0398_),
    .Y(_0442_),
    .A1(net571),
    .A2(_0346_));
 sg13g2_nor2b_1 _4069_ (.A(_0442_),
    .B_N(_0441_),
    .Y(_0443_));
 sg13g2_nand2_1 _4070_ (.Y(_0444_),
    .A(net622),
    .B(_0912_));
 sg13g2_o21ai_1 _4071_ (.B1(_0444_),
    .Y(_0445_),
    .A1(_0912_),
    .A2(_0334_));
 sg13g2_mux2_1 _4072_ (.A0(net631),
    .A1(_0360_),
    .S(_0945_),
    .X(_0446_));
 sg13g2_nand2_1 _4073_ (.Y(_0447_),
    .A(net635),
    .B(_0736_));
 sg13g2_nand3_1 _4074_ (.B(_2647_),
    .C(_0221_),
    .A(_2668_),
    .Y(_0448_));
 sg13g2_a21oi_1 _4075_ (.A1(_0747_),
    .A2(_1438_),
    .Y(_0449_),
    .B1(_0226_));
 sg13g2_or2_1 _4076_ (.X(_0451_),
    .B(_0449_),
    .A(_0448_));
 sg13g2_a21oi_1 _4077_ (.A1(_0447_),
    .A2(_0451_),
    .Y(_0452_),
    .B1(_0446_));
 sg13g2_a21oi_1 _4078_ (.A1(net627),
    .A2(net547),
    .Y(_0453_),
    .B1(_0452_));
 sg13g2_xnor2_1 _4079_ (.Y(_0454_),
    .A(_0445_),
    .B(_0453_));
 sg13g2_nand3_1 _4080_ (.B(_0447_),
    .C(_0451_),
    .A(_0446_),
    .Y(_0455_));
 sg13g2_nand2b_1 _4081_ (.Y(_0456_),
    .B(_0455_),
    .A_N(_0452_));
 sg13g2_nor2_1 _4082_ (.A(net588),
    .B(_0456_),
    .Y(_0457_));
 sg13g2_xnor2_1 _4083_ (.Y(_0458_),
    .A(_0448_),
    .B(_0449_));
 sg13g2_nor2_1 _4084_ (.A(net592),
    .B(_0458_),
    .Y(_0459_));
 sg13g2_and2_1 _4085_ (.A(_2647_),
    .B(_2682_),
    .X(_0460_));
 sg13g2_xnor2_1 _4086_ (.Y(_0462_),
    .A(net558),
    .B(_0460_));
 sg13g2_a221oi_1 _4087_ (.B2(_2682_),
    .C1(_0423_),
    .B1(_0703_),
    .A1(net559),
    .Y(_0463_),
    .A2(_0692_));
 sg13g2_a221oi_1 _4088_ (.B2(net595),
    .C1(_0463_),
    .B1(_0462_),
    .A1(_1021_),
    .Y(_0464_),
    .A2(_0425_));
 sg13g2_nor2_1 _4089_ (.A(net595),
    .B(_0462_),
    .Y(_0465_));
 sg13g2_nor3_1 _4090_ (.A(_0459_),
    .B(_0464_),
    .C(_0465_),
    .Y(_0466_));
 sg13g2_a21oi_1 _4091_ (.A1(net592),
    .A2(_0458_),
    .Y(_0467_),
    .B1(_0466_));
 sg13g2_a22oi_1 _4092_ (.Y(_0468_),
    .B1(_0456_),
    .B2(net589),
    .A2(_0454_),
    .A1(net584));
 sg13g2_o21ai_1 _4093_ (.B1(_0468_),
    .Y(_0469_),
    .A1(_0457_),
    .A2(_0467_));
 sg13g2_o21ai_1 _4094_ (.B1(_0469_),
    .Y(_0470_),
    .A1(net585),
    .A2(_0454_));
 sg13g2_o21ai_1 _4095_ (.B1(_0444_),
    .Y(_0471_),
    .A1(_0445_),
    .A2(_0453_));
 sg13g2_nor2_1 _4096_ (.A(net629),
    .B(_0659_),
    .Y(_0473_));
 sg13g2_a21oi_1 _4097_ (.A1(_1744_),
    .A2(_0235_),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_xnor2_1 _4098_ (.Y(_0475_),
    .A(_0471_),
    .B(_0474_));
 sg13g2_nand2_1 _4099_ (.Y(_0476_),
    .A(net581),
    .B(_0475_));
 sg13g2_a21oi_1 _4100_ (.A1(_0471_),
    .A2(_0474_),
    .Y(_0477_),
    .B1(_0473_));
 sg13g2_xnor2_1 _4101_ (.Y(_0478_),
    .A(net613),
    .B(_1723_));
 sg13g2_nor2_1 _4102_ (.A(_0477_),
    .B(_0478_),
    .Y(_0479_));
 sg13g2_xnor2_1 _4103_ (.Y(_0480_),
    .A(_0477_),
    .B(_0478_));
 sg13g2_nor2_1 _4104_ (.A(net581),
    .B(_0475_),
    .Y(_0481_));
 sg13g2_o21ai_1 _4105_ (.B1(_0476_),
    .Y(_0482_),
    .A1(_0470_),
    .A2(_0481_));
 sg13g2_o21ai_1 _4106_ (.B1(_0482_),
    .Y(_0484_),
    .A1(net575),
    .A2(_0480_));
 sg13g2_xor2_1 _4107_ (.B(net607),
    .A(net617),
    .X(_0485_));
 sg13g2_a21oi_1 _4108_ (.A1(net613),
    .A2(_1723_),
    .Y(_0486_),
    .B1(_0479_));
 sg13g2_xnor2_1 _4109_ (.Y(_0487_),
    .A(_0485_),
    .B(_0486_));
 sg13g2_a22oi_1 _4110_ (.Y(_0488_),
    .B1(_0487_),
    .B2(net571),
    .A2(_0480_),
    .A1(net575));
 sg13g2_a21oi_1 _4111_ (.A1(net555),
    .A2(_0479_),
    .Y(_0489_),
    .B1(net608));
 sg13g2_mux2_1 _4112_ (.A0(_0604_),
    .A1(net612),
    .S(_0489_),
    .X(_0490_));
 sg13g2_o21ai_1 _4113_ (.B1(_0490_),
    .Y(_0491_),
    .A1(net571),
    .A2(_0487_));
 sg13g2_a21oi_1 _4114_ (.A1(_0484_),
    .A2(_0488_),
    .Y(_0492_),
    .B1(_0491_));
 sg13g2_nor2_2 _4115_ (.A(_0443_),
    .B(_0492_),
    .Y(_0493_));
 sg13g2_xnor2_1 _4116_ (.Y(_0495_),
    .A(net538),
    .B(_0493_));
 sg13g2_nor3_1 _4117_ (.A(_2577_),
    .B(net473),
    .C(_0495_),
    .Y(_0496_));
 sg13g2_inv_1 _4118_ (.Y(_0497_),
    .A(_0496_));
 sg13g2_nor2b_2 _4119_ (.A(_0065_),
    .B_N(_0098_),
    .Y(_0498_));
 sg13g2_nand2b_1 _4120_ (.Y(_0499_),
    .B(_0098_),
    .A_N(net550));
 sg13g2_nor2_1 _4121_ (.A(_0307_),
    .B(net471),
    .Y(_0500_));
 sg13g2_a22oi_1 _4122_ (.Y(_0501_),
    .B1(_2420_),
    .B2(net533),
    .A2(net502),
    .A1(_2646_));
 sg13g2_nand2_2 _4123_ (.Y(_0502_),
    .A(_1251_),
    .B(net498));
 sg13g2_and2_1 _4124_ (.A(_1284_),
    .B(_0502_),
    .X(_0503_));
 sg13g2_o21ai_1 _4125_ (.B1(_0501_),
    .Y(_0504_),
    .A1(net509),
    .A2(_0503_));
 sg13g2_nand2_1 _4126_ (.Y(_0506_),
    .A(_2027_),
    .B(_0502_));
 sg13g2_xnor2_1 _4127_ (.Y(_0507_),
    .A(_2027_),
    .B(_0502_));
 sg13g2_a22oi_1 _4128_ (.Y(_0508_),
    .B1(_0507_),
    .B2(net512),
    .A2(_0503_),
    .A1(net509));
 sg13g2_or2_1 _4129_ (.X(_0509_),
    .B(_0506_),
    .A(net503));
 sg13g2_xnor2_1 _4130_ (.Y(_0510_),
    .A(net504),
    .B(_0506_));
 sg13g2_nor2_1 _4131_ (.A(net510),
    .B(_0510_),
    .Y(_0511_));
 sg13g2_a21oi_1 _4132_ (.A1(_0504_),
    .A2(_0508_),
    .Y(_0512_),
    .B1(_0511_));
 sg13g2_o21ai_1 _4133_ (.B1(_0512_),
    .Y(_0513_),
    .A1(net512),
    .A2(_0507_));
 sg13g2_nand2_1 _4134_ (.Y(_0514_),
    .A(net462),
    .B(_0509_));
 sg13g2_xnor2_1 _4135_ (.Y(_0515_),
    .A(net462),
    .B(_0509_));
 sg13g2_o21ai_1 _4136_ (.B1(_0513_),
    .Y(_0517_),
    .A1(net514),
    .A2(_0515_));
 sg13g2_a21oi_1 _4137_ (.A1(net510),
    .A2(_0510_),
    .Y(_0518_),
    .B1(_0517_));
 sg13g2_nor2_1 _4138_ (.A(_1581_),
    .B(_0514_),
    .Y(_0519_));
 sg13g2_xnor2_1 _4139_ (.Y(_0520_),
    .A(_1581_),
    .B(_0514_));
 sg13g2_a221oi_1 _4140_ (.B2(net508),
    .C1(_0518_),
    .B1(_0520_),
    .A1(net514),
    .Y(_0521_),
    .A2(_0515_));
 sg13g2_nor2_1 _4141_ (.A(net508),
    .B(_0520_),
    .Y(_0522_));
 sg13g2_xnor2_1 _4142_ (.Y(_0523_),
    .A(net461),
    .B(_0519_));
 sg13g2_a21oi_1 _4143_ (.A1(_0989_),
    .A2(_0523_),
    .Y(_0524_),
    .B1(_0522_));
 sg13g2_nand2_1 _4144_ (.Y(_0525_),
    .A(_0331_),
    .B(_0524_));
 sg13g2_a21oi_1 _4145_ (.A1(_0703_),
    .A2(net513),
    .Y(_0526_),
    .B1(_2635_));
 sg13g2_nor2_1 _4146_ (.A(_0714_),
    .B(_0526_),
    .Y(_0528_));
 sg13g2_nand2_1 _4147_ (.Y(_0529_),
    .A(net638),
    .B(_0714_));
 sg13g2_nand2_1 _4148_ (.Y(_0530_),
    .A(net510),
    .B(_0529_));
 sg13g2_nand2_1 _4149_ (.Y(_0531_),
    .A(_0758_),
    .B(_0530_));
 sg13g2_nand2_1 _4150_ (.Y(_0532_),
    .A(_1897_),
    .B(_0531_));
 sg13g2_a21oi_1 _4151_ (.A1(net510),
    .A2(_0529_),
    .Y(_0533_),
    .B1(net515));
 sg13g2_xnor2_1 _4152_ (.Y(_0534_),
    .A(net514),
    .B(_0530_));
 sg13g2_o21ai_1 _4153_ (.B1(_0528_),
    .Y(_0535_),
    .A1(_1897_),
    .A2(_0531_));
 sg13g2_a22oi_1 _4154_ (.Y(_0536_),
    .B1(_0535_),
    .B2(_0532_),
    .A2(_0534_),
    .A1(net502));
 sg13g2_nor2_1 _4155_ (.A(net502),
    .B(_0534_),
    .Y(_0537_));
 sg13g2_nand2_1 _4156_ (.Y(_0539_),
    .A(net508),
    .B(_0533_));
 sg13g2_xnor2_1 _4157_ (.Y(_0540_),
    .A(net508),
    .B(_0533_));
 sg13g2_nor2_1 _4158_ (.A(net499),
    .B(_0540_),
    .Y(_0541_));
 sg13g2_nor3_1 _4159_ (.A(_0536_),
    .B(_0537_),
    .C(_0541_),
    .Y(_0542_));
 sg13g2_xnor2_1 _4160_ (.Y(_0543_),
    .A(_0978_),
    .B(_0539_));
 sg13g2_a221oi_1 _4161_ (.B2(net506),
    .C1(_0542_),
    .B1(_0543_),
    .A1(net499),
    .Y(_0544_),
    .A2(_0540_));
 sg13g2_nand2b_1 _4162_ (.Y(_0545_),
    .B(_0539_),
    .A_N(_2105_));
 sg13g2_a21o_1 _4163_ (.A2(_0539_),
    .A1(_0989_),
    .B1(net461),
    .X(_0546_));
 sg13g2_and2_1 _4164_ (.A(_0545_),
    .B(_0546_),
    .X(_0547_));
 sg13g2_or2_1 _4165_ (.X(_0548_),
    .B(_0547_),
    .A(net503));
 sg13g2_o21ai_1 _4166_ (.B1(_0548_),
    .Y(_0550_),
    .A1(net506),
    .A2(_0543_));
 sg13g2_nor2_1 _4167_ (.A(_0626_),
    .B(_1734_),
    .Y(_0551_));
 sg13g2_o21ai_1 _4168_ (.B1(_0258_),
    .Y(_0552_),
    .A1(_0967_),
    .A2(_0551_));
 sg13g2_nor2_1 _4169_ (.A(net621),
    .B(_0615_),
    .Y(_0553_));
 sg13g2_nand2_1 _4170_ (.Y(_0554_),
    .A(_0670_),
    .B(_0552_));
 sg13g2_o21ai_1 _4171_ (.B1(_1570_),
    .Y(_0555_),
    .A1(_0545_),
    .A2(_0554_));
 sg13g2_nand2_1 _4172_ (.Y(_0556_),
    .A(_0545_),
    .B(_0554_));
 sg13g2_a21o_1 _4173_ (.A2(_0556_),
    .A1(_1581_),
    .B1(net462),
    .X(_0557_));
 sg13g2_a21oi_1 _4174_ (.A1(_2533_),
    .A2(_0556_),
    .Y(_0558_),
    .B1(_0555_));
 sg13g2_a221oi_1 _4175_ (.B2(_0557_),
    .C1(_0558_),
    .B1(_0555_),
    .A1(net503),
    .Y(_0559_),
    .A2(_0547_));
 sg13g2_o21ai_1 _4176_ (.B1(_0559_),
    .Y(_0561_),
    .A1(_0544_),
    .A2(_0550_));
 sg13g2_o21ai_1 _4177_ (.B1(_0561_),
    .Y(_0562_),
    .A1(_0521_),
    .A2(_0525_));
 sg13g2_nand3_1 _4178_ (.B(_1240_),
    .C(_2112_),
    .A(net593),
    .Y(_0563_));
 sg13g2_o21ai_1 _4179_ (.B1(_0563_),
    .Y(_0564_),
    .A1(_0615_),
    .A2(_0529_));
 sg13g2_nor3_1 _4180_ (.A(_0519_),
    .B(_0556_),
    .C(_0564_),
    .Y(_0565_));
 sg13g2_nand2_2 _4181_ (.Y(_0566_),
    .A(_0562_),
    .B(_0565_));
 sg13g2_nor3_1 _4182_ (.A(_0307_),
    .B(net471),
    .C(_0566_),
    .Y(_0567_));
 sg13g2_nand3_1 _4183_ (.B(net578),
    .C(net593),
    .A(net573),
    .Y(_0568_));
 sg13g2_and4_1 _4184_ (.A(net563),
    .B(_0549_),
    .C(_1152_),
    .D(_0568_),
    .X(_0569_));
 sg13g2_nand4_1 _4185_ (.B(_0549_),
    .C(_1152_),
    .A(net564),
    .Y(_0570_),
    .D(_0568_));
 sg13g2_or3_1 _4186_ (.A(net557),
    .B(net476),
    .C(_0310_),
    .X(_0572_));
 sg13g2_a221oi_1 _4187_ (.B2(_0311_),
    .C1(_0309_),
    .B1(_0308_),
    .A1(net621),
    .Y(_0573_),
    .A2(_0240_));
 sg13g2_a221oi_1 _4188_ (.B2(_0573_),
    .C1(_0250_),
    .B1(_0572_),
    .A1(net556),
    .Y(_0574_),
    .A2(net475));
 sg13g2_nor2_2 _4189_ (.A(_0253_),
    .B(_0574_),
    .Y(_0575_));
 sg13g2_inv_1 _4190_ (.Y(_0576_),
    .A(_0575_));
 sg13g2_nor3_1 _4191_ (.A(_0340_),
    .B(net495),
    .C(_0575_),
    .Y(_0577_));
 sg13g2_nor2_2 _4192_ (.A(_1548_),
    .B(_2572_),
    .Y(_0578_));
 sg13g2_nand2b_2 _4193_ (.Y(_0579_),
    .B(_1537_),
    .A_N(_2572_));
 sg13g2_nor2_2 _4194_ (.A(net539),
    .B(_0578_),
    .Y(_0580_));
 sg13g2_nand2_2 _4195_ (.Y(_0581_),
    .A(net548),
    .B(net468));
 sg13g2_and2_1 _4196_ (.A(net588),
    .B(net594),
    .X(_0583_));
 sg13g2_nand2_1 _4197_ (.Y(_0584_),
    .A(net590),
    .B(net594));
 sg13g2_a21oi_1 _4198_ (.A1(_1537_),
    .A2(_0583_),
    .Y(_0585_),
    .B1(_0581_));
 sg13g2_and4_1 _4199_ (.A(_0219_),
    .B(_2565_),
    .C(_0576_),
    .D(_0585_),
    .X(_0586_));
 sg13g2_nor2_1 _4200_ (.A(_0450_),
    .B(net471),
    .Y(_0587_));
 sg13g2_a21o_1 _4201_ (.A2(_0500_),
    .A1(_0681_),
    .B1(_0587_),
    .X(_0588_));
 sg13g2_nand2_2 _4202_ (.Y(_0589_),
    .A(_0296_),
    .B(_2625_));
 sg13g2_nand3_1 _4203_ (.B(_2625_),
    .C(_0498_),
    .A(_0175_),
    .Y(_0590_));
 sg13g2_a21oi_1 _4204_ (.A1(_2626_),
    .A2(net457),
    .Y(_0591_),
    .B1(net470));
 sg13g2_nor2_1 _4205_ (.A(_2569_),
    .B(net577),
    .Y(_0592_));
 sg13g2_nand2_1 _4206_ (.Y(_0594_),
    .A(net544),
    .B(_0592_));
 sg13g2_o21ai_1 _4207_ (.B1(net593),
    .Y(_0595_),
    .A1(net596),
    .A2(_0425_));
 sg13g2_o21ai_1 _4208_ (.B1(_2573_),
    .Y(_0596_),
    .A1(_0594_),
    .A2(_0595_));
 sg13g2_nand2_1 _4209_ (.Y(_0597_),
    .A(net590),
    .B(net599));
 sg13g2_a21oi_1 _4210_ (.A1(_0584_),
    .A2(_0597_),
    .Y(_0598_),
    .B1(_1262_));
 sg13g2_a21oi_1 _4211_ (.A1(net577),
    .A2(_0598_),
    .Y(_0599_),
    .B1(_2605_));
 sg13g2_nor2_2 _4212_ (.A(net563),
    .B(_0599_),
    .Y(_0600_));
 sg13g2_nand2b_2 _4213_ (.Y(_0601_),
    .B(net568),
    .A_N(_0599_));
 sg13g2_and2_1 _4214_ (.A(net566),
    .B(_0596_),
    .X(_0602_));
 sg13g2_nand2_2 _4215_ (.Y(_0603_),
    .A(net566),
    .B(_0596_));
 sg13g2_nand2_2 _4216_ (.Y(_0605_),
    .A(_0600_),
    .B(net447));
 sg13g2_nand2_2 _4217_ (.Y(_0606_),
    .A(net563),
    .B(_2587_));
 sg13g2_nor2_1 _4218_ (.A(net590),
    .B(_1273_),
    .Y(_0607_));
 sg13g2_o21ai_1 _4219_ (.B1(net579),
    .Y(_0608_),
    .A1(_1273_),
    .A2(net544));
 sg13g2_nand2_2 _4220_ (.Y(_0609_),
    .A(net541),
    .B(_0608_));
 sg13g2_and2_1 _4221_ (.A(net541),
    .B(_0608_),
    .X(_0610_));
 sg13g2_nand3_1 _4222_ (.B(net593),
    .C(_1251_),
    .A(net572),
    .Y(_0611_));
 sg13g2_o21ai_1 _4223_ (.B1(net572),
    .Y(_0612_),
    .A1(net579),
    .A2(net544));
 sg13g2_and3_2 _4224_ (.X(_0613_),
    .A(net562),
    .B(_0611_),
    .C(_0612_));
 sg13g2_nand3_1 _4225_ (.B(_0611_),
    .C(_0612_),
    .A(net562),
    .Y(_0614_));
 sg13g2_nand2_2 _4226_ (.Y(_0616_),
    .A(net454),
    .B(net467));
 sg13g2_and2_1 _4227_ (.A(_0605_),
    .B(_0616_),
    .X(_0617_));
 sg13g2_a21oi_1 _4228_ (.A1(net538),
    .A2(_0588_),
    .Y(_0618_),
    .B1(_0567_));
 sg13g2_a221oi_1 _4229_ (.B2(_0617_),
    .C1(_0586_),
    .B1(_0591_),
    .A1(_0569_),
    .Y(_0619_),
    .A2(_0577_));
 sg13g2_nand2_2 _4230_ (.Y(_0620_),
    .A(_0362_),
    .B(_0264_));
 sg13g2_nor2_2 _4231_ (.A(_2019_),
    .B(_0583_),
    .Y(_0621_));
 sg13g2_nor2_1 _4232_ (.A(net637),
    .B(_2329_),
    .Y(_0622_));
 sg13g2_nand2b_1 _4233_ (.Y(_0623_),
    .B(_0305_),
    .A_N(_0622_));
 sg13g2_o21ai_1 _4234_ (.B1(_0623_),
    .Y(_0624_),
    .A1(_2679_),
    .A2(net497));
 sg13g2_o21ai_1 _4235_ (.B1(_0624_),
    .Y(_0625_),
    .A1(net633),
    .A2(_0621_));
 sg13g2_nand2_1 _4236_ (.Y(_0627_),
    .A(net498),
    .B(_0312_));
 sg13g2_o21ai_1 _4237_ (.B1(_0627_),
    .Y(_0628_),
    .A1(net585),
    .A2(net498));
 sg13g2_a22oi_1 _4238_ (.Y(_0629_),
    .B1(_0628_),
    .B2(net626),
    .A2(_0621_),
    .A1(net633));
 sg13g2_a21oi_1 _4239_ (.A1(net475),
    .A2(_0271_),
    .Y(_0630_),
    .B1(_0289_));
 sg13g2_or2_1 _4240_ (.X(_0631_),
    .B(_0628_),
    .A(net626));
 sg13g2_o21ai_1 _4241_ (.B1(_0631_),
    .Y(_0632_),
    .A1(net624),
    .A2(_0630_));
 sg13g2_a21oi_1 _4242_ (.A1(_0625_),
    .A2(_0629_),
    .Y(_0633_),
    .B1(_0632_));
 sg13g2_o21ai_1 _4243_ (.B1(_0245_),
    .Y(_0634_),
    .A1(_2329_),
    .A2(_0288_));
 sg13g2_xnor2_1 _4244_ (.Y(_0635_),
    .A(_0246_),
    .B(_0289_));
 sg13g2_a221oi_1 _4245_ (.B2(net616),
    .C1(_0633_),
    .B1(_0635_),
    .A1(net621),
    .Y(_0636_),
    .A2(_0630_));
 sg13g2_nand2b_1 _4246_ (.Y(_0638_),
    .B(net552),
    .A_N(_0634_));
 sg13g2_o21ai_1 _4247_ (.B1(_0638_),
    .Y(_0639_),
    .A1(net616),
    .A2(_0635_));
 sg13g2_a21oi_1 _4248_ (.A1(net614),
    .A2(_0634_),
    .Y(_0640_),
    .B1(net606));
 sg13g2_o21ai_1 _4249_ (.B1(_0640_),
    .Y(_0641_),
    .A1(_0636_),
    .A2(_0639_));
 sg13g2_nand2_1 _4250_ (.Y(_0642_),
    .A(net534),
    .B(_0641_));
 sg13g2_a21oi_1 _4251_ (.A1(_0255_),
    .A2(_0642_),
    .Y(_0643_),
    .B1(_0620_));
 sg13g2_nand2_1 _4252_ (.Y(_0644_),
    .A(_2583_),
    .B(_2606_));
 sg13g2_nor2_2 _4253_ (.A(_0340_),
    .B(net471),
    .Y(_0645_));
 sg13g2_a21oi_2 _4254_ (.B1(_2606_),
    .Y(_0646_),
    .A2(net493),
    .A1(net546));
 sg13g2_inv_1 _4255_ (.Y(_0647_),
    .A(_0646_));
 sg13g2_nor2_2 _4256_ (.A(net539),
    .B(_2606_),
    .Y(_0649_));
 sg13g2_nand2_2 _4257_ (.Y(_0650_),
    .A(net549),
    .B(net522));
 sg13g2_o21ai_1 _4258_ (.B1(net549),
    .Y(_0651_),
    .A1(net492),
    .A2(net468));
 sg13g2_o21ai_1 _4259_ (.B1(_0645_),
    .Y(_0652_),
    .A1(_0647_),
    .A2(_0651_));
 sg13g2_nor2b_1 _4260_ (.A(_0652_),
    .B_N(_0644_),
    .Y(_0653_));
 sg13g2_nand2_1 _4261_ (.Y(_0654_),
    .A(_0516_),
    .B(_0583_));
 sg13g2_o21ai_1 _4262_ (.B1(net541),
    .Y(_0655_),
    .A1(_0527_),
    .A2(_0584_));
 sg13g2_a21oi_1 _4263_ (.A1(_0516_),
    .A2(_0583_),
    .Y(_0656_),
    .B1(_2604_));
 sg13g2_nor3_1 _4264_ (.A(_0527_),
    .B(_1548_),
    .C(_2019_),
    .Y(_0657_));
 sg13g2_nor2_2 _4265_ (.A(net539),
    .B(_0657_),
    .Y(_0658_));
 sg13g2_or2_1 _4266_ (.X(_0660_),
    .B(_0657_),
    .A(net539));
 sg13g2_nor2_2 _4267_ (.A(net535),
    .B(net451),
    .Y(_0661_));
 sg13g2_inv_1 _4268_ (.Y(_0662_),
    .A(_0661_));
 sg13g2_nand2_2 _4269_ (.Y(_0663_),
    .A(_0252_),
    .B(_2567_));
 sg13g2_nor2_2 _4270_ (.A(net471),
    .B(_0663_),
    .Y(_0664_));
 sg13g2_o21ai_1 _4271_ (.B1(_0664_),
    .Y(_0665_),
    .A1(net520),
    .A2(_0661_));
 sg13g2_nand2_2 _4272_ (.Y(_0666_),
    .A(_0208_),
    .B(_2625_));
 sg13g2_nor2_2 _4273_ (.A(net477),
    .B(_0666_),
    .Y(_0667_));
 sg13g2_nand2_2 _4274_ (.Y(_0668_),
    .A(_0252_),
    .B(_2625_));
 sg13g2_nor3_2 _4275_ (.A(net528),
    .B(net477),
    .C(_0668_),
    .Y(_0669_));
 sg13g2_a21oi_1 _4276_ (.A1(net535),
    .A2(_0667_),
    .Y(_0671_),
    .B1(_0669_));
 sg13g2_nand2_1 _4277_ (.Y(_0672_),
    .A(_0665_),
    .B(_0671_));
 sg13g2_and2_1 _4278_ (.A(net550),
    .B(_0417_),
    .X(_0673_));
 sg13g2_nand2_1 _4279_ (.Y(_0674_),
    .A(net550),
    .B(_0417_));
 sg13g2_nor2_2 _4280_ (.A(_0666_),
    .B(net465),
    .Y(_0675_));
 sg13g2_nor2_2 _4281_ (.A(_0267_),
    .B(net465),
    .Y(_0676_));
 sg13g2_nor2_1 _4282_ (.A(_0274_),
    .B(net478),
    .Y(_0677_));
 sg13g2_nor3_1 _4283_ (.A(_0675_),
    .B(_0676_),
    .C(_0677_),
    .Y(_0678_));
 sg13g2_nand2_2 _4284_ (.Y(_0679_),
    .A(_0263_),
    .B(_0296_));
 sg13g2_nor2_2 _4285_ (.A(net473),
    .B(_0679_),
    .Y(_0680_));
 sg13g2_nand2_2 _4286_ (.Y(_0682_),
    .A(_0362_),
    .B(_0673_));
 sg13g2_o21ai_1 _4287_ (.B1(_0678_),
    .Y(_0683_),
    .A1(net526),
    .A2(_0682_));
 sg13g2_a21o_1 _4288_ (.A2(_0680_),
    .A1(_0649_),
    .B1(_0683_),
    .X(_0684_));
 sg13g2_nor3_1 _4289_ (.A(_0653_),
    .B(_0672_),
    .C(_0684_),
    .Y(_0685_));
 sg13g2_a21oi_2 _4290_ (.B1(_0569_),
    .Y(_0686_),
    .A2(_2036_),
    .A1(_2033_));
 sg13g2_a21o_2 _4291_ (.A2(_2036_),
    .A1(_2033_),
    .B1(_0569_),
    .X(_0687_));
 sg13g2_nor2_2 _4292_ (.A(net479),
    .B(_0267_),
    .Y(_0688_));
 sg13g2_nand3_1 _4293_ (.B(net450),
    .C(_0688_),
    .A(net455),
    .Y(_0689_));
 sg13g2_nand2_1 _4294_ (.Y(_0690_),
    .A(net447),
    .B(net450));
 sg13g2_nand2_2 _4295_ (.Y(_0691_),
    .A(_0208_),
    .B(_2567_));
 sg13g2_nor2_1 _4296_ (.A(net469),
    .B(_0691_),
    .Y(_0693_));
 sg13g2_nand3_1 _4297_ (.B(_2567_),
    .C(_0498_),
    .A(_0208_),
    .Y(_0694_));
 sg13g2_nand3_1 _4298_ (.B(_0690_),
    .C(_0693_),
    .A(_0616_),
    .Y(_0695_));
 sg13g2_nor2_2 _4299_ (.A(net457),
    .B(net465),
    .Y(_0696_));
 sg13g2_inv_1 _4300_ (.Y(_0697_),
    .A(_0696_));
 sg13g2_o21ai_1 _4301_ (.B1(net485),
    .Y(_0698_),
    .A1(net519),
    .A2(_0661_));
 sg13g2_nor2_2 _4302_ (.A(net565),
    .B(_0612_),
    .Y(_0699_));
 sg13g2_nand2_1 _4303_ (.Y(_0700_),
    .A(_2583_),
    .B(_0699_));
 sg13g2_a21oi_1 _4304_ (.A1(net524),
    .A2(_0700_),
    .Y(_0701_),
    .B1(net534));
 sg13g2_nor4_1 _4305_ (.A(net516),
    .B(_0340_),
    .C(net531),
    .D(_0701_),
    .Y(_0702_));
 sg13g2_a21oi_1 _4306_ (.A1(_0696_),
    .A2(_0698_),
    .Y(_0704_),
    .B1(_0702_));
 sg13g2_nand4_1 _4307_ (.B(_0689_),
    .C(_0695_),
    .A(_0685_),
    .Y(_0705_),
    .D(_0704_));
 sg13g2_nor2_2 _4308_ (.A(net495),
    .B(_2626_),
    .Y(_0706_));
 sg13g2_nor2_1 _4309_ (.A(net480),
    .B(_0602_),
    .Y(_0707_));
 sg13g2_nor2_2 _4310_ (.A(_0600_),
    .B(net452),
    .Y(_0708_));
 sg13g2_nand2_2 _4311_ (.Y(_0709_),
    .A(net487),
    .B(net452));
 sg13g2_o21ai_1 _4312_ (.B1(_0706_),
    .Y(_0710_),
    .A1(_0707_),
    .A2(_0708_));
 sg13g2_nand2_1 _4313_ (.Y(_0711_),
    .A(_1537_),
    .B(_2572_));
 sg13g2_o21ai_1 _4314_ (.B1(net590),
    .Y(_0712_),
    .A1(net599),
    .A2(_1273_));
 sg13g2_o21ai_1 _4315_ (.B1(_0580_),
    .Y(_0713_),
    .A1(_0711_),
    .A2(_0712_));
 sg13g2_inv_1 _4316_ (.Y(_0715_),
    .A(net446));
 sg13g2_nor2_2 _4317_ (.A(_0687_),
    .B(net446),
    .Y(_0716_));
 sg13g2_nand2_1 _4318_ (.Y(_0717_),
    .A(net450),
    .B(_0715_));
 sg13g2_nand2_2 _4319_ (.Y(_0718_),
    .A(net447),
    .B(net454));
 sg13g2_nor2_1 _4320_ (.A(_0716_),
    .B(net444),
    .Y(_0719_));
 sg13g2_or2_1 _4321_ (.X(_0720_),
    .B(net444),
    .A(_0716_));
 sg13g2_nor2_1 _4322_ (.A(_2577_),
    .B(net469),
    .Y(_0721_));
 sg13g2_nand2_1 _4323_ (.Y(_0722_),
    .A(_0720_),
    .B(_0721_));
 sg13g2_nand2_1 _4324_ (.Y(_0723_),
    .A(net583),
    .B(_0592_));
 sg13g2_a21oi_1 _4325_ (.A1(_2591_),
    .A2(_0595_),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_nor3_1 _4326_ (.A(net563),
    .B(_1141_),
    .C(_1262_),
    .Y(_0726_));
 sg13g2_nor2_1 _4327_ (.A(net525),
    .B(_0726_),
    .Y(_0727_));
 sg13g2_o21ai_1 _4328_ (.B1(_0727_),
    .Y(_0728_),
    .A1(net532),
    .A2(_0724_));
 sg13g2_nor2_1 _4329_ (.A(net495),
    .B(_0663_),
    .Y(_0729_));
 sg13g2_nor3_1 _4330_ (.A(net495),
    .B(_0613_),
    .C(_0663_),
    .Y(_0730_));
 sg13g2_nand2_1 _4331_ (.Y(_0731_),
    .A(_0728_),
    .B(_0730_));
 sg13g2_nor2_1 _4332_ (.A(net546),
    .B(_0578_),
    .Y(_0732_));
 sg13g2_o21ai_1 _4333_ (.B1(net522),
    .Y(_0733_),
    .A1(net546),
    .A2(_0578_));
 sg13g2_nor2_1 _4334_ (.A(net495),
    .B(_0691_),
    .Y(_0734_));
 sg13g2_a22oi_1 _4335_ (.Y(_0735_),
    .B1(_0733_),
    .B2(_0734_),
    .A2(_0730_),
    .A1(_0728_));
 sg13g2_nand3_1 _4336_ (.B(_0722_),
    .C(_0735_),
    .A(_0710_),
    .Y(_0737_));
 sg13g2_nor2_1 _4337_ (.A(_0705_),
    .B(_0737_),
    .Y(_0738_));
 sg13g2_nor2_2 _4338_ (.A(_2577_),
    .B(net477),
    .Y(_0739_));
 sg13g2_nand2_2 _4339_ (.Y(_0740_),
    .A(_2576_),
    .B(_2627_));
 sg13g2_nor2_2 _4340_ (.A(_0230_),
    .B(net479),
    .Y(_0741_));
 sg13g2_nor2_2 _4341_ (.A(_0340_),
    .B(_2628_),
    .Y(_0742_));
 sg13g2_a22oi_1 _4342_ (.Y(_0743_),
    .B1(_0742_),
    .B2(_0662_),
    .A2(_0741_),
    .A1(_0658_));
 sg13g2_a22oi_1 _4343_ (.Y(_0744_),
    .B1(_0740_),
    .B2(_0743_),
    .A2(net519),
    .A1(net480));
 sg13g2_nor2_1 _4344_ (.A(net478),
    .B(_0663_),
    .Y(_0745_));
 sg13g2_nor2_2 _4345_ (.A(net545),
    .B(_0581_),
    .Y(_0746_));
 sg13g2_nand2_2 _4346_ (.Y(_0748_),
    .A(net532),
    .B(_0580_));
 sg13g2_nor2_2 _4347_ (.A(_2568_),
    .B(net478),
    .Y(_0749_));
 sg13g2_nand2_1 _4348_ (.Y(_0750_),
    .A(net483),
    .B(_0699_));
 sg13g2_nor2_1 _4349_ (.A(net526),
    .B(net491),
    .Y(_0751_));
 sg13g2_nand2_2 _4350_ (.Y(_0752_),
    .A(net531),
    .B(net483));
 sg13g2_a21o_2 _4351_ (.A2(net544),
    .A1(net580),
    .B1(_2604_),
    .X(_0753_));
 sg13g2_a21oi_2 _4352_ (.B1(_2604_),
    .Y(_0754_),
    .A2(net544),
    .A1(net580));
 sg13g2_nand3_1 _4353_ (.B(_0752_),
    .C(_0753_),
    .A(_0750_),
    .Y(_0755_));
 sg13g2_a22oi_1 _4354_ (.Y(_0756_),
    .B1(_0749_),
    .B2(_0755_),
    .A2(net445),
    .A1(_0745_));
 sg13g2_nand2_2 _4355_ (.Y(_0757_),
    .A(_2643_),
    .B(_2647_));
 sg13g2_nand3_1 _4356_ (.B(_2552_),
    .C(_0757_),
    .A(_0923_),
    .Y(_0759_));
 sg13g2_a21oi_1 _4357_ (.A1(net629),
    .A2(_2552_),
    .Y(_0760_),
    .B1(net609));
 sg13g2_nand2_1 _4358_ (.Y(_0761_),
    .A(_0759_),
    .B(_0760_));
 sg13g2_nand3_1 _4359_ (.B(_0759_),
    .C(_0760_),
    .A(net553),
    .Y(_0762_));
 sg13g2_inv_1 _4360_ (.Y(_0763_),
    .A(_0762_));
 sg13g2_nor2_2 _4361_ (.A(net472),
    .B(_0668_),
    .Y(_0764_));
 sg13g2_a22oi_1 _4362_ (.Y(_0765_),
    .B1(_0763_),
    .B2(_0764_),
    .A2(net447),
    .A1(_0318_));
 sg13g2_nand2_1 _4363_ (.Y(_0766_),
    .A(_0756_),
    .B(_0765_));
 sg13g2_nor2_1 _4364_ (.A(net455),
    .B(_0707_),
    .Y(_0767_));
 sg13g2_nor2_2 _4365_ (.A(net482),
    .B(_0614_),
    .Y(_0768_));
 sg13g2_nor2_2 _4366_ (.A(net452),
    .B(_0768_),
    .Y(_0770_));
 sg13g2_o21ai_1 _4367_ (.B1(net454),
    .Y(_0771_),
    .A1(net480),
    .A2(_0614_));
 sg13g2_nor2_2 _4368_ (.A(_0373_),
    .B(net477),
    .Y(_0772_));
 sg13g2_nand2_2 _4369_ (.Y(_0773_),
    .A(_0362_),
    .B(_2627_));
 sg13g2_nor3_1 _4370_ (.A(_0767_),
    .B(_0771_),
    .C(_0773_),
    .Y(_0774_));
 sg13g2_nand2_2 _4371_ (.Y(_0775_),
    .A(net488),
    .B(_0602_));
 sg13g2_nor2_1 _4372_ (.A(_0373_),
    .B(net469),
    .Y(_0776_));
 sg13g2_nand3_1 _4373_ (.B(_0775_),
    .C(_0776_),
    .A(net453),
    .Y(_0777_));
 sg13g2_a21oi_1 _4374_ (.A1(net487),
    .A2(_0716_),
    .Y(_0778_),
    .B1(_0777_));
 sg13g2_nor4_1 _4375_ (.A(_0744_),
    .B(_0766_),
    .C(_0774_),
    .D(_0778_),
    .Y(_0779_));
 sg13g2_nor2_2 _4376_ (.A(_0373_),
    .B(net496),
    .Y(_0781_));
 sg13g2_nand2_1 _4377_ (.Y(_0782_),
    .A(_0362_),
    .B(_2565_));
 sg13g2_nor2_1 _4378_ (.A(net548),
    .B(net489),
    .Y(_0783_));
 sg13g2_nor2_1 _4379_ (.A(net545),
    .B(_0783_),
    .Y(_0784_));
 sg13g2_inv_1 _4380_ (.Y(_0785_),
    .A(_0784_));
 sg13g2_nand2_1 _4381_ (.Y(_0786_),
    .A(_0781_),
    .B(_0785_));
 sg13g2_nor2_2 _4382_ (.A(net472),
    .B(net457),
    .Y(_0787_));
 sg13g2_a22oi_1 _4383_ (.Y(_0788_),
    .B1(_0787_),
    .B2(net548),
    .A2(_0785_),
    .A1(_0781_));
 sg13g2_nand3_1 _4384_ (.B(_0263_),
    .C(_2565_),
    .A(_0252_),
    .Y(_0789_));
 sg13g2_nor2_1 _4385_ (.A(net538),
    .B(_0789_),
    .Y(_0790_));
 sg13g2_nor2_2 _4386_ (.A(_2626_),
    .B(net473),
    .Y(_0792_));
 sg13g2_o21ai_1 _4387_ (.B1(_0792_),
    .Y(_0793_),
    .A1(net481),
    .A2(_0733_));
 sg13g2_nand3b_1 _4388_ (.B(_0793_),
    .C(_0788_),
    .Y(_0794_),
    .A_N(_0790_));
 sg13g2_nor2_2 _4389_ (.A(net496),
    .B(net457),
    .Y(_0795_));
 sg13g2_nor4_1 _4390_ (.A(net539),
    .B(net495),
    .C(_2608_),
    .D(net457),
    .Y(_0796_));
 sg13g2_nand2_2 _4391_ (.Y(_0797_),
    .A(_0266_),
    .B(_0498_));
 sg13g2_nor3_1 _4392_ (.A(_0578_),
    .B(_0783_),
    .C(_0797_),
    .Y(_0798_));
 sg13g2_nand2_2 _4393_ (.Y(_0799_),
    .A(_0219_),
    .B(_0498_));
 sg13g2_nor2_2 _4394_ (.A(net479),
    .B(_0691_),
    .Y(_0800_));
 sg13g2_nand2_1 _4395_ (.Y(_0801_),
    .A(net445),
    .B(_0800_));
 sg13g2_o21ai_1 _4396_ (.B1(_0801_),
    .Y(_0803_),
    .A1(_0748_),
    .A2(_0799_));
 sg13g2_nor4_1 _4397_ (.A(_0794_),
    .B(_0796_),
    .C(_0798_),
    .D(_0803_),
    .Y(_0804_));
 sg13g2_nand3_1 _4398_ (.B(_0439_),
    .C(_2627_),
    .A(_0153_),
    .Y(_0805_));
 sg13g2_nand2_2 _4399_ (.Y(_0806_),
    .A(net534),
    .B(net491));
 sg13g2_nand2_1 _4400_ (.Y(_0807_),
    .A(net521),
    .B(_0806_));
 sg13g2_nand2_1 _4401_ (.Y(_0808_),
    .A(net489),
    .B(net519));
 sg13g2_a21o_1 _4402_ (.A2(_0808_),
    .A1(_0807_),
    .B1(_0805_),
    .X(_0809_));
 sg13g2_nor2_2 _4403_ (.A(net478),
    .B(_0589_),
    .Y(_0810_));
 sg13g2_nor2_2 _4404_ (.A(_2577_),
    .B(net465),
    .Y(_0811_));
 sg13g2_a22oi_1 _4405_ (.Y(_0812_),
    .B1(_0811_),
    .B2(net523),
    .A2(_0810_),
    .A1(net546));
 sg13g2_nor2_2 _4406_ (.A(_0340_),
    .B(net472),
    .Y(_0814_));
 sg13g2_nor4_1 _4407_ (.A(net477),
    .B(_0580_),
    .C(net457),
    .D(_0783_),
    .Y(_0815_));
 sg13g2_a21oi_1 _4408_ (.A1(net534),
    .A2(_0814_),
    .Y(_0816_),
    .B1(_0815_));
 sg13g2_nand4_1 _4409_ (.B(_0809_),
    .C(_0812_),
    .A(_0804_),
    .Y(_0817_),
    .D(_0816_));
 sg13g2_nor2_1 _4410_ (.A(net496),
    .B(_0267_),
    .Y(_0818_));
 sg13g2_nand2_2 _4411_ (.Y(_0819_),
    .A(_2565_),
    .B(_0266_));
 sg13g2_nor2_2 _4412_ (.A(_1185_),
    .B(net492),
    .Y(_0820_));
 sg13g2_nor3_1 _4413_ (.A(_2574_),
    .B(_0699_),
    .C(_0820_),
    .Y(_0821_));
 sg13g2_nor2_1 _4414_ (.A(_0274_),
    .B(net472),
    .Y(_0822_));
 sg13g2_a21oi_2 _4415_ (.B1(_2580_),
    .Y(_0823_),
    .A2(_2447_),
    .A1(_2591_));
 sg13g2_a21oi_2 _4416_ (.B1(net525),
    .Y(_0825_),
    .A2(_0823_),
    .A1(net568));
 sg13g2_nand3_1 _4417_ (.B(_0822_),
    .C(_0825_),
    .A(net521),
    .Y(_0826_));
 sg13g2_o21ai_1 _4418_ (.B1(_0826_),
    .Y(_0827_),
    .A1(_0819_),
    .A2(_0821_));
 sg13g2_nor2_2 _4419_ (.A(_0274_),
    .B(net465),
    .Y(_0828_));
 sg13g2_nor2_2 _4420_ (.A(net478),
    .B(_0679_),
    .Y(_0829_));
 sg13g2_o21ai_1 _4421_ (.B1(net548),
    .Y(_0830_),
    .A1(_0828_),
    .A2(_0829_));
 sg13g2_nor2_2 _4422_ (.A(net496),
    .B(_0668_),
    .Y(_0831_));
 sg13g2_o21ai_1 _4423_ (.B1(net570),
    .Y(_0832_),
    .A1(net490),
    .A2(_0581_));
 sg13g2_a21oi_1 _4424_ (.A1(net532),
    .A2(net482),
    .Y(_0833_),
    .B1(net570));
 sg13g2_nand2_1 _4425_ (.Y(_0834_),
    .A(_0549_),
    .B(_0833_));
 sg13g2_nand2_1 _4426_ (.Y(_0836_),
    .A(_0832_),
    .B(_0834_));
 sg13g2_nand2_1 _4427_ (.Y(_0837_),
    .A(_0831_),
    .B(_0836_));
 sg13g2_o21ai_1 _4428_ (.B1(_0837_),
    .Y(_0838_),
    .A1(net546),
    .A2(_0830_));
 sg13g2_nor2_2 _4429_ (.A(net474),
    .B(_0691_),
    .Y(_0839_));
 sg13g2_o21ai_1 _4430_ (.B1(_0733_),
    .Y(_0840_),
    .A1(net483),
    .A2(_0650_));
 sg13g2_inv_1 _4431_ (.Y(_0841_),
    .A(_0840_));
 sg13g2_nor2_2 _4432_ (.A(_2626_),
    .B(net465),
    .Y(_0842_));
 sg13g2_a22oi_1 _4433_ (.Y(_0843_),
    .B1(_0841_),
    .B2(_0842_),
    .A2(_0839_),
    .A1(_0651_));
 sg13g2_nor2_2 _4434_ (.A(_0230_),
    .B(net473),
    .Y(_0844_));
 sg13g2_nand2_2 _4435_ (.Y(_0845_),
    .A(_0687_),
    .B(_0844_));
 sg13g2_nor2_1 _4436_ (.A(_0663_),
    .B(net465),
    .Y(_0847_));
 sg13g2_nand3_1 _4437_ (.B(_2567_),
    .C(_0673_),
    .A(_0252_),
    .Y(_0848_));
 sg13g2_nand2_1 _4438_ (.Y(_0849_),
    .A(_0840_),
    .B(_0847_));
 sg13g2_nor2_2 _4439_ (.A(net496),
    .B(_0679_),
    .Y(_0850_));
 sg13g2_nor2_2 _4440_ (.A(net474),
    .B(_0666_),
    .Y(_0851_));
 sg13g2_or2_1 _4441_ (.X(_0852_),
    .B(_0851_),
    .A(_0850_));
 sg13g2_a21oi_1 _4442_ (.A1(net493),
    .A2(net525),
    .Y(_0853_),
    .B1(net531));
 sg13g2_nor2_2 _4443_ (.A(net531),
    .B(net524),
    .Y(_0854_));
 sg13g2_nand2_2 _4444_ (.Y(_0855_),
    .A(net527),
    .B(net542));
 sg13g2_a21oi_1 _4445_ (.A1(_0752_),
    .A2(_0855_),
    .Y(_0856_),
    .B1(_0395_));
 sg13g2_nand2_2 _4446_ (.Y(_0858_),
    .A(net545),
    .B(_2605_));
 sg13g2_nor2_1 _4447_ (.A(net473),
    .B(_0663_),
    .Y(_0859_));
 sg13g2_or2_1 _4448_ (.X(_0860_),
    .B(_0663_),
    .A(net474));
 sg13g2_a221oi_1 _4449_ (.B2(_0859_),
    .C1(_0856_),
    .B1(_0858_),
    .A1(_0852_),
    .Y(_0861_),
    .A2(_0853_));
 sg13g2_nand4_1 _4450_ (.B(_0845_),
    .C(_0849_),
    .A(_0843_),
    .Y(_0862_),
    .D(_0861_));
 sg13g2_nor4_1 _4451_ (.A(_0817_),
    .B(_0827_),
    .C(_0838_),
    .D(_0862_),
    .Y(_0863_));
 sg13g2_and2_1 _4452_ (.A(_0605_),
    .B(net446),
    .X(_0864_));
 sg13g2_nor2_2 _4453_ (.A(_0687_),
    .B(_0864_),
    .Y(_0865_));
 sg13g2_nor3_1 _4454_ (.A(net480),
    .B(net467),
    .C(_0865_),
    .Y(_0866_));
 sg13g2_nor2_1 _4455_ (.A(_0307_),
    .B(net477),
    .Y(_0867_));
 sg13g2_nor4_1 _4456_ (.A(_0307_),
    .B(net477),
    .C(net452),
    .D(_0866_),
    .Y(_0869_));
 sg13g2_nor2_2 _4457_ (.A(_0274_),
    .B(net470),
    .Y(_0870_));
 sg13g2_o21ai_1 _4458_ (.B1(_0864_),
    .Y(_0871_),
    .A1(net487),
    .A2(_0602_));
 sg13g2_nand2_1 _4459_ (.Y(_0872_),
    .A(_2584_),
    .B(_0687_));
 sg13g2_nand2_1 _4460_ (.Y(_0873_),
    .A(net487),
    .B(_0687_));
 sg13g2_nand3_1 _4461_ (.B(_0871_),
    .C(_0873_),
    .A(net454),
    .Y(_0874_));
 sg13g2_nand2_2 _4462_ (.Y(_0875_),
    .A(net480),
    .B(_0610_));
 sg13g2_nand3_1 _4463_ (.B(_0874_),
    .C(_0875_),
    .A(_0616_),
    .Y(_0876_));
 sg13g2_a21oi_1 _4464_ (.A1(_0870_),
    .A2(_0876_),
    .Y(_0877_),
    .B1(_0869_));
 sg13g2_nand4_1 _4465_ (.B(_0779_),
    .C(_0863_),
    .A(_0738_),
    .Y(_0878_),
    .D(_0877_));
 sg13g2_nand4_1 _4466_ (.B(net455),
    .C(net447),
    .A(net480),
    .Y(_0880_),
    .D(net450));
 sg13g2_o21ai_1 _4467_ (.B1(_0600_),
    .Y(_0881_),
    .A1(net487),
    .A2(_0602_));
 sg13g2_nand4_1 _4468_ (.B(_0770_),
    .C(_0880_),
    .A(_0717_),
    .Y(_0882_),
    .D(_0881_));
 sg13g2_nand2_1 _4469_ (.Y(_0883_),
    .A(_0461_),
    .B(_0709_));
 sg13g2_nor2b_1 _4470_ (.A(_0883_),
    .B_N(_0882_),
    .Y(_0884_));
 sg13g2_nor2_1 _4471_ (.A(net469),
    .B(_0668_),
    .Y(_0885_));
 sg13g2_nand2_1 _4472_ (.Y(_0886_),
    .A(_0616_),
    .B(_0885_));
 sg13g2_o21ai_1 _4473_ (.B1(net637),
    .Y(_0887_),
    .A1(net646),
    .A2(net642));
 sg13g2_nand2_2 _4474_ (.Y(_0888_),
    .A(net557),
    .B(_0887_));
 sg13g2_nand3_1 _4475_ (.B(_0333_),
    .C(_0888_),
    .A(_0331_),
    .Y(_0889_));
 sg13g2_nand3_1 _4476_ (.B(_0359_),
    .C(_0757_),
    .A(_1734_),
    .Y(_0891_));
 sg13g2_nor3_1 _4477_ (.A(net552),
    .B(net606),
    .C(_2582_),
    .Y(_0892_));
 sg13g2_nand3_1 _4478_ (.B(_2636_),
    .C(_0891_),
    .A(net554),
    .Y(_0893_));
 sg13g2_a21oi_1 _4479_ (.A1(_0681_),
    .A2(_0889_),
    .Y(_0894_),
    .B1(_0893_));
 sg13g2_nand3_1 _4480_ (.B(net490),
    .C(_0889_),
    .A(_0681_),
    .Y(_0895_));
 sg13g2_a221oi_1 _4481_ (.B2(_0894_),
    .C1(_0716_),
    .B1(_0892_),
    .A1(_1755_),
    .Y(_0896_),
    .A2(_2584_));
 sg13g2_nand4_1 _4482_ (.B(_0762_),
    .C(_0895_),
    .A(net456),
    .Y(_0897_),
    .D(_0896_));
 sg13g2_a21oi_1 _4483_ (.A1(_0605_),
    .A2(_0897_),
    .Y(_0898_),
    .B1(net452));
 sg13g2_nor2_1 _4484_ (.A(_0886_),
    .B(_0898_),
    .Y(_0899_));
 sg13g2_nor2_1 _4485_ (.A(net495),
    .B(_0666_),
    .Y(_0900_));
 sg13g2_nand3_1 _4486_ (.B(_2565_),
    .C(_2625_),
    .A(_0208_),
    .Y(_0902_));
 sg13g2_nor2_1 _4487_ (.A(net452),
    .B(_0902_),
    .Y(_0903_));
 sg13g2_nand2b_2 _4488_ (.Y(_0904_),
    .B(_0264_),
    .A_N(_2568_));
 sg13g2_nor3_2 _4489_ (.A(_0600_),
    .B(net467),
    .C(_0904_),
    .Y(_0905_));
 sg13g2_a22oi_1 _4490_ (.Y(_0906_),
    .B1(_0905_),
    .B2(_0717_),
    .A2(_0903_),
    .A1(_0605_));
 sg13g2_a21o_1 _4491_ (.A2(net467),
    .A1(net482),
    .B1(_0906_),
    .X(_0907_));
 sg13g2_nor2_1 _4492_ (.A(_2568_),
    .B(net466),
    .Y(_0908_));
 sg13g2_nand3_1 _4493_ (.B(_2567_),
    .C(_0673_),
    .A(_0296_),
    .Y(_0909_));
 sg13g2_nor2_2 _4494_ (.A(_0340_),
    .B(net466),
    .Y(_0910_));
 sg13g2_a21oi_2 _4495_ (.B1(net590),
    .Y(_0911_),
    .A2(_1207_),
    .A1(net594));
 sg13g2_o21ai_1 _4496_ (.B1(_0580_),
    .Y(_0913_),
    .A1(_0711_),
    .A2(_0911_));
 sg13g2_inv_1 _4497_ (.Y(_0914_),
    .A(_0913_));
 sg13g2_nor2_2 _4498_ (.A(_0307_),
    .B(net472),
    .Y(_0915_));
 sg13g2_nor2b_2 _4499_ (.A(_0913_),
    .B_N(_0915_),
    .Y(_0916_));
 sg13g2_nor2_2 _4500_ (.A(_0450_),
    .B(net473),
    .Y(_0917_));
 sg13g2_inv_1 _4501_ (.Y(_0918_),
    .A(_0917_));
 sg13g2_nand2_1 _4502_ (.Y(_0919_),
    .A(net534),
    .B(_0917_));
 sg13g2_nand2_2 _4503_ (.Y(_0920_),
    .A(_0219_),
    .B(_0673_));
 sg13g2_inv_1 _4504_ (.Y(_0921_),
    .A(_0920_));
 sg13g2_nor2_1 _4505_ (.A(net523),
    .B(_0920_),
    .Y(_0922_));
 sg13g2_o21ai_1 _4506_ (.B1(_0919_),
    .Y(_0924_),
    .A1(_0718_),
    .A2(_0909_));
 sg13g2_nor4_2 _4507_ (.A(_0910_),
    .B(_0916_),
    .C(_0922_),
    .Y(_0925_),
    .D(_0924_));
 sg13g2_nor2_2 _4508_ (.A(net470),
    .B(_0666_),
    .Y(_0926_));
 sg13g2_a22oi_1 _4509_ (.Y(_0927_),
    .B1(net446),
    .B2(net447),
    .A2(net467),
    .A1(net453));
 sg13g2_nor2_1 _4510_ (.A(_2568_),
    .B(net469),
    .Y(_0928_));
 sg13g2_nand2_1 _4511_ (.Y(_0929_),
    .A(_0720_),
    .B(_0928_));
 sg13g2_a22oi_1 _4512_ (.Y(_0930_),
    .B1(_0928_),
    .B2(_0720_),
    .A2(_0927_),
    .A1(_0926_));
 sg13g2_o21ai_1 _4513_ (.B1(_0505_),
    .Y(_0931_),
    .A1(_0607_),
    .A2(_0723_));
 sg13g2_nand2_1 _4514_ (.Y(_0932_),
    .A(net568),
    .B(_0931_));
 sg13g2_o21ai_1 _4515_ (.B1(_0505_),
    .Y(_0933_),
    .A1(_0911_),
    .A2(_0932_));
 sg13g2_nand2_1 _4516_ (.Y(_0935_),
    .A(net560),
    .B(_2036_));
 sg13g2_a21oi_1 _4517_ (.A1(_2032_),
    .A2(_0935_),
    .Y(_0936_),
    .B1(_1109_));
 sg13g2_a21oi_1 _4518_ (.A1(_0913_),
    .A2(_0933_),
    .Y(_0937_),
    .B1(_0936_));
 sg13g2_nor2_1 _4519_ (.A(net530),
    .B(_0937_),
    .Y(_0938_));
 sg13g2_a21oi_1 _4520_ (.A1(net541),
    .A2(_0911_),
    .Y(_0939_),
    .B1(_2606_));
 sg13g2_inv_1 _4521_ (.Y(_0940_),
    .A(_0939_));
 sg13g2_nor3_1 _4522_ (.A(net466),
    .B(_0691_),
    .C(_0938_),
    .Y(_0941_));
 sg13g2_nor2_2 _4523_ (.A(_0668_),
    .B(net466),
    .Y(_0942_));
 sg13g2_o21ai_1 _4524_ (.B1(net446),
    .Y(_0943_),
    .A1(net653),
    .A2(_0600_));
 sg13g2_nand4_1 _4525_ (.B(_0614_),
    .C(_0872_),
    .A(net482),
    .Y(_0944_),
    .D(_0943_));
 sg13g2_nand2b_1 _4526_ (.Y(_0946_),
    .B(_0944_),
    .A_N(net444));
 sg13g2_a22oi_1 _4527_ (.Y(_0947_),
    .B1(_0942_),
    .B2(_0946_),
    .A2(_0941_),
    .A1(_0939_));
 sg13g2_nand4_1 _4528_ (.B(_0925_),
    .C(_0930_),
    .A(_0907_),
    .Y(_0948_),
    .D(_0947_));
 sg13g2_nor4_2 _4529_ (.A(_0878_),
    .B(_0884_),
    .C(_0899_),
    .Y(_0949_),
    .D(_0948_));
 sg13g2_a21oi_1 _4530_ (.A1(net562),
    .A2(_2573_),
    .Y(_0950_),
    .B1(_2613_));
 sg13g2_xnor2_1 _4531_ (.Y(_0951_),
    .A(_2613_),
    .B(net529));
 sg13g2_nor2_1 _4532_ (.A(net560),
    .B(net529),
    .Y(_0952_));
 sg13g2_xnor2_1 _4533_ (.Y(_0953_),
    .A(net560),
    .B(net529));
 sg13g2_a22oi_1 _4534_ (.Y(_0954_),
    .B1(_0953_),
    .B2(net638),
    .A2(_0951_),
    .A1(net642));
 sg13g2_nand2b_1 _4535_ (.Y(_0955_),
    .B(_2690_),
    .A_N(_0951_));
 sg13g2_xnor2_1 _4536_ (.Y(_0957_),
    .A(_2624_),
    .B(net529));
 sg13g2_nor2_1 _4537_ (.A(net646),
    .B(_0957_),
    .Y(_0958_));
 sg13g2_xnor2_1 _4538_ (.Y(_0959_),
    .A(net603),
    .B(net529));
 sg13g2_nand2_1 _4539_ (.Y(_0960_),
    .A(net559),
    .B(_0959_));
 sg13g2_a21oi_1 _4540_ (.A1(net646),
    .A2(_0957_),
    .Y(_0961_),
    .B1(_0960_));
 sg13g2_nor2_1 _4541_ (.A(_0958_),
    .B(_0961_),
    .Y(_0962_));
 sg13g2_nand2_1 _4542_ (.Y(_0963_),
    .A(_0955_),
    .B(_0962_));
 sg13g2_xnor2_1 _4543_ (.Y(_0964_),
    .A(_2591_),
    .B(net529));
 sg13g2_nor2_1 _4544_ (.A(net636),
    .B(_0953_),
    .Y(_0965_));
 sg13g2_a21oi_1 _4545_ (.A1(_0954_),
    .A2(_0963_),
    .Y(_0966_),
    .B1(_0965_));
 sg13g2_o21ai_1 _4546_ (.B1(_0966_),
    .Y(_0968_),
    .A1(net633),
    .A2(_0964_));
 sg13g2_nand2_1 _4547_ (.Y(_0969_),
    .A(net583),
    .B(_2604_));
 sg13g2_nor2_1 _4548_ (.A(net583),
    .B(net545),
    .Y(_0970_));
 sg13g2_inv_1 _4549_ (.Y(_0971_),
    .A(_0970_));
 sg13g2_o21ai_1 _4550_ (.B1(_0971_),
    .Y(_0972_),
    .A1(_2580_),
    .A2(_2604_));
 sg13g2_a22oi_1 _4551_ (.Y(_0973_),
    .B1(_0972_),
    .B2(net627),
    .A2(_0964_),
    .A1(net634));
 sg13g2_xnor2_1 _4552_ (.Y(_0974_),
    .A(net528),
    .B(_0238_));
 sg13g2_xnor2_1 _4553_ (.Y(_0975_),
    .A(net530),
    .B(_0238_));
 sg13g2_nor2_1 _4554_ (.A(net627),
    .B(_0972_),
    .Y(_0976_));
 sg13g2_a221oi_1 _4555_ (.B2(net556),
    .C1(_0976_),
    .B1(_0975_),
    .A1(_0968_),
    .Y(_0977_),
    .A2(_0973_));
 sg13g2_a221oi_1 _4556_ (.B2(net621),
    .C1(_0977_),
    .B1(_0974_),
    .A1(net616),
    .Y(_0979_),
    .A2(_0244_));
 sg13g2_a22oi_1 _4557_ (.Y(_0980_),
    .B1(_0593_),
    .B2(_1109_),
    .A2(_0527_),
    .A1(_2569_));
 sg13g2_o21ai_1 _4558_ (.B1(_2605_),
    .Y(_0981_),
    .A1(_0582_),
    .A2(_1098_));
 sg13g2_nand2_1 _4559_ (.Y(_0982_),
    .A(net552),
    .B(_0980_));
 sg13g2_o21ai_1 _4560_ (.B1(_0982_),
    .Y(_0983_),
    .A1(net619),
    .A2(_0244_));
 sg13g2_nor2_1 _4561_ (.A(_0979_),
    .B(_0983_),
    .Y(_0984_));
 sg13g2_a21oi_1 _4562_ (.A1(net614),
    .A2(_0981_),
    .Y(_0985_),
    .B1(net606));
 sg13g2_nor2b_1 _4563_ (.A(_0984_),
    .B_N(_0985_),
    .Y(_0986_));
 sg13g2_inv_2 _4564_ (.Y(_0987_),
    .A(_0986_));
 sg13g2_nor2_2 _4565_ (.A(_0450_),
    .B(net465),
    .Y(_0988_));
 sg13g2_nor2_2 _4566_ (.A(_0307_),
    .B(net466),
    .Y(_0990_));
 sg13g2_a21oi_1 _4567_ (.A1(_0854_),
    .A2(_0988_),
    .Y(_0991_),
    .B1(_0990_));
 sg13g2_a21oi_1 _4568_ (.A1(_0855_),
    .A2(_0987_),
    .Y(_0992_),
    .B1(_0991_));
 sg13g2_nand3_1 _4569_ (.B(_0619_),
    .C(_0949_),
    .A(_0618_),
    .Y(_0993_));
 sg13g2_nor4_1 _4570_ (.A(_0496_),
    .B(_0643_),
    .C(_0992_),
    .D(_0993_),
    .Y(_0994_));
 sg13g2_and3_1 _4571_ (.X(_0995_),
    .A(_0327_),
    .B(_0422_),
    .C(_0994_));
 sg13g2_nand4_1 _4572_ (.B(_2616_),
    .C(_2631_),
    .A(_2593_),
    .Y(_0996_),
    .D(_0995_));
 sg13g2_nor2b_2 _4573_ (.A(_0637_),
    .B_N(_0996_),
    .Y(uo_out[4]));
 sg13g2_o21ai_1 _4574_ (.B1(net570),
    .Y(_0997_),
    .A1(_1273_),
    .A2(net544));
 sg13g2_nand3_1 _4575_ (.B(_2607_),
    .C(_0997_),
    .A(net542),
    .Y(_0998_));
 sg13g2_a21oi_1 _4576_ (.A1(_2600_),
    .A2(_0998_),
    .Y(_1000_),
    .B1(_2601_));
 sg13g2_o21ai_1 _4577_ (.B1(_1000_),
    .Y(_1001_),
    .A1(_2599_),
    .A2(_2611_));
 sg13g2_o21ai_1 _4578_ (.B1(net538),
    .Y(_1002_),
    .A1(net565),
    .A2(_0612_));
 sg13g2_nand3b_1 _4579_ (.B(_0641_),
    .C(_1002_),
    .Y(_1003_),
    .A_N(_0325_));
 sg13g2_nor2_2 _4580_ (.A(net497),
    .B(_2421_),
    .Y(_1004_));
 sg13g2_xnor2_1 _4581_ (.Y(_1005_),
    .A(_0225_),
    .B(_1004_));
 sg13g2_nor2_1 _4582_ (.A(net633),
    .B(_1005_),
    .Y(_1006_));
 sg13g2_a21oi_1 _4583_ (.A1(_2679_),
    .A2(_2448_),
    .Y(_1007_),
    .B1(_0279_));
 sg13g2_a21oi_1 _4584_ (.A1(net637),
    .A2(_2449_),
    .Y(_1008_),
    .B1(_1007_));
 sg13g2_nand2b_2 _4585_ (.Y(_1009_),
    .B(_0270_),
    .A_N(_1004_));
 sg13g2_o21ai_1 _4586_ (.B1(net585),
    .Y(_1011_),
    .A1(_0224_),
    .A2(_1004_));
 sg13g2_and2_1 _4587_ (.A(_1009_),
    .B(_1011_),
    .X(_1012_));
 sg13g2_a22oi_1 _4588_ (.Y(_1013_),
    .B1(_1012_),
    .B2(net626),
    .A2(_1005_),
    .A1(net634));
 sg13g2_o21ai_1 _4589_ (.B1(_1013_),
    .Y(_1014_),
    .A1(_1006_),
    .A2(_1008_));
 sg13g2_xnor2_1 _4590_ (.Y(_1015_),
    .A(net475),
    .B(_1009_));
 sg13g2_nor2_1 _4591_ (.A(net622),
    .B(_1015_),
    .Y(_1016_));
 sg13g2_nor2_1 _4592_ (.A(net628),
    .B(_1012_),
    .Y(_1017_));
 sg13g2_nor2_1 _4593_ (.A(_1016_),
    .B(_1017_),
    .Y(_1018_));
 sg13g2_a21oi_1 _4594_ (.A1(net475),
    .A2(_1009_),
    .Y(_1019_),
    .B1(_0245_));
 sg13g2_nand3_1 _4595_ (.B(_0245_),
    .C(_1009_),
    .A(net475),
    .Y(_1020_));
 sg13g2_nor2b_1 _4596_ (.A(_1019_),
    .B_N(_1020_),
    .Y(_1022_));
 sg13g2_and2_1 _4597_ (.A(net617),
    .B(_1022_),
    .X(_1023_));
 sg13g2_a221oi_1 _4598_ (.B2(_1014_),
    .C1(_1023_),
    .B1(_1018_),
    .A1(net622),
    .Y(_1024_),
    .A2(_1015_));
 sg13g2_nor2_1 _4599_ (.A(net617),
    .B(_1022_),
    .Y(_1025_));
 sg13g2_nor2_1 _4600_ (.A(net611),
    .B(_1019_),
    .Y(_1026_));
 sg13g2_nor3_1 _4601_ (.A(_1024_),
    .B(_1025_),
    .C(_1026_),
    .Y(_1027_));
 sg13g2_a21oi_1 _4602_ (.A1(net611),
    .A2(_1019_),
    .Y(_1028_),
    .B1(net607));
 sg13g2_nor2b_1 _4603_ (.A(_1027_),
    .B_N(_1028_),
    .Y(_1029_));
 sg13g2_a21oi_1 _4604_ (.A1(_0641_),
    .A2(_1029_),
    .Y(_1030_),
    .B1(_0575_));
 sg13g2_and2_1 _4605_ (.A(_0300_),
    .B(_1030_),
    .X(_1031_));
 sg13g2_a21oi_1 _4606_ (.A1(_1003_),
    .A2(_1031_),
    .Y(_1033_),
    .B1(_0269_));
 sg13g2_nand3_1 _4607_ (.B(_0770_),
    .C(_0881_),
    .A(_0461_),
    .Y(_1034_));
 sg13g2_nor2_1 _4608_ (.A(_0645_),
    .B(_0839_),
    .Y(_1035_));
 sg13g2_a21oi_2 _4609_ (.B1(_0606_),
    .Y(_1036_),
    .A2(_2446_),
    .A1(_1131_));
 sg13g2_nor2_1 _4610_ (.A(_0825_),
    .B(_0931_),
    .Y(_1037_));
 sg13g2_nor4_1 _4611_ (.A(_0274_),
    .B(net472),
    .C(_1036_),
    .D(_1037_),
    .Y(_1038_));
 sg13g2_o21ai_1 _4612_ (.B1(_1002_),
    .Y(_1039_),
    .A1(_0814_),
    .A2(_0818_));
 sg13g2_or2_1 _4613_ (.X(_1040_),
    .B(_0867_),
    .A(_0776_));
 sg13g2_a21oi_1 _4614_ (.A1(_0913_),
    .A2(_0933_),
    .Y(_1041_),
    .B1(net530));
 sg13g2_a21oi_1 _4615_ (.A1(net560),
    .A2(_2036_),
    .Y(_1042_),
    .B1(_1141_));
 sg13g2_nor2_2 _4616_ (.A(_0606_),
    .B(_1042_),
    .Y(_1044_));
 sg13g2_nor3_2 _4617_ (.A(net466),
    .B(_0691_),
    .C(_1044_),
    .Y(_1045_));
 sg13g2_o21ai_1 _4618_ (.B1(_1045_),
    .Y(_1046_),
    .A1(_0940_),
    .A2(_1041_));
 sg13g2_nand2_1 _4619_ (.Y(_1047_),
    .A(_0662_),
    .B(_0739_));
 sg13g2_nand3_1 _4620_ (.B(_0805_),
    .C(_1047_),
    .A(_0743_),
    .Y(_1048_));
 sg13g2_o21ai_1 _4621_ (.B1(net453),
    .Y(_1049_),
    .A1(net467),
    .A2(_0865_));
 sg13g2_nor3_1 _4622_ (.A(_2568_),
    .B(net469),
    .C(_1049_),
    .Y(_1050_));
 sg13g2_a21oi_1 _4623_ (.A1(_0590_),
    .A2(_0904_),
    .Y(_1051_),
    .B1(net444));
 sg13g2_and3_1 _4624_ (.X(_1052_),
    .A(net456),
    .B(_0728_),
    .C(_0729_));
 sg13g2_nor2_2 _4625_ (.A(net520),
    .B(net451),
    .Y(_1053_));
 sg13g2_nand2_2 _4626_ (.Y(_1055_),
    .A(net521),
    .B(_0658_));
 sg13g2_nor3_1 _4627_ (.A(_2577_),
    .B(net472),
    .C(_1055_),
    .Y(_1056_));
 sg13g2_a21o_1 _4628_ (.A2(_0734_),
    .A1(_0649_),
    .B1(_1056_),
    .X(_1057_));
 sg13g2_nor3_1 _4629_ (.A(_1051_),
    .B(_1052_),
    .C(_1057_),
    .Y(_1058_));
 sg13g2_nand2b_1 _4630_ (.Y(_1059_),
    .B(net453),
    .A_N(_0864_));
 sg13g2_nor2_1 _4631_ (.A(_0694_),
    .B(_1059_),
    .Y(_1060_));
 sg13g2_o21ai_1 _4632_ (.B1(_0831_),
    .Y(_1061_),
    .A1(net530),
    .A2(_0834_));
 sg13g2_nor2_2 _4633_ (.A(_0650_),
    .B(_0799_),
    .Y(_1062_));
 sg13g2_a21oi_1 _4634_ (.A1(net539),
    .A2(net492),
    .Y(_1063_),
    .B1(_0797_));
 sg13g2_nor2_1 _4635_ (.A(net446),
    .B(_0773_),
    .Y(_1064_));
 sg13g2_nand2_1 _4636_ (.Y(_1066_),
    .A(net455),
    .B(_0870_));
 sg13g2_nand4_1 _4637_ (.B(_0750_),
    .C(_0752_),
    .A(_0749_),
    .Y(_1067_),
    .D(_0753_));
 sg13g2_nand2_1 _4638_ (.Y(_1068_),
    .A(_0395_),
    .B(_2578_));
 sg13g2_a21oi_1 _4639_ (.A1(net445),
    .A2(_0800_),
    .Y(_1069_),
    .B1(_0669_));
 sg13g2_nor2_2 _4640_ (.A(_0450_),
    .B(net496),
    .Y(_1070_));
 sg13g2_nor2_2 _4641_ (.A(net466),
    .B(_0679_),
    .Y(_1071_));
 sg13g2_nor3_1 _4642_ (.A(_0721_),
    .B(_0885_),
    .C(_0926_),
    .Y(_1072_));
 sg13g2_or2_1 _4643_ (.X(_1073_),
    .B(_1072_),
    .A(net444));
 sg13g2_nor2_1 _4644_ (.A(net481),
    .B(net468),
    .Y(_1074_));
 sg13g2_nor4_2 _4645_ (.A(net539),
    .B(net477),
    .C(_0663_),
    .Y(_1075_),
    .D(_1074_));
 sg13g2_nor2_2 _4646_ (.A(net471),
    .B(_0679_),
    .Y(_1077_));
 sg13g2_nor3_1 _4647_ (.A(_0781_),
    .B(_0787_),
    .C(_1077_),
    .Y(_1078_));
 sg13g2_nor2_1 _4648_ (.A(_2594_),
    .B(_0234_),
    .Y(_1079_));
 sg13g2_nand2_1 _4649_ (.Y(_1080_),
    .A(_0888_),
    .B(_1079_));
 sg13g2_and2_1 _4650_ (.A(_2596_),
    .B(_1080_),
    .X(_1081_));
 sg13g2_nand2_2 _4651_ (.Y(_1082_),
    .A(_2596_),
    .B(_1080_));
 sg13g2_o21ai_1 _4652_ (.B1(_1073_),
    .Y(_1083_),
    .A1(_0581_),
    .A2(_1078_));
 sg13g2_a22oi_1 _4653_ (.Y(_1084_),
    .B1(_1075_),
    .B2(net532),
    .A2(_1068_),
    .A1(net542));
 sg13g2_nand3_1 _4654_ (.B(_1067_),
    .C(_1084_),
    .A(_0925_),
    .Y(_1085_));
 sg13g2_a221oi_1 _4655_ (.B2(_0285_),
    .C1(_1063_),
    .B1(net464),
    .A1(_0785_),
    .Y(_1086_),
    .A2(_0810_));
 sg13g2_o21ai_1 _4656_ (.B1(_1086_),
    .Y(_1088_),
    .A1(_2606_),
    .A2(_0860_));
 sg13g2_a22oi_1 _4657_ (.Y(_1089_),
    .B1(_0855_),
    .B2(_0811_),
    .A2(_0828_),
    .A1(_0649_));
 sg13g2_o21ai_1 _4658_ (.B1(_1089_),
    .Y(_1090_),
    .A1(_0918_),
    .A2(_0932_));
 sg13g2_nor4_1 _4659_ (.A(_0684_),
    .B(_1085_),
    .C(_1088_),
    .D(_1090_),
    .Y(_1091_));
 sg13g2_a22oi_1 _4660_ (.Y(_1092_),
    .B1(_1048_),
    .B2(_0808_),
    .A2(_0944_),
    .A1(_0942_));
 sg13g2_a22oi_1 _4661_ (.Y(_1093_),
    .B1(_0915_),
    .B2(_0933_),
    .A2(_0844_),
    .A1(_0690_));
 sg13g2_o21ai_1 _4662_ (.B1(_1061_),
    .Y(_1094_),
    .A1(_0651_),
    .A2(_1035_));
 sg13g2_a21oi_1 _4663_ (.A1(_0688_),
    .A2(_0716_),
    .Y(_1095_),
    .B1(_1094_));
 sg13g2_nand2b_1 _4664_ (.Y(_1096_),
    .B(_0789_),
    .A_N(_0667_));
 sg13g2_a22oi_1 _4665_ (.Y(_1097_),
    .B1(_1096_),
    .B2(_0658_),
    .A2(_1040_),
    .A1(_0614_));
 sg13g2_a21oi_1 _4666_ (.A1(net447),
    .A2(_0900_),
    .Y(_1099_),
    .B1(_1038_));
 sg13g2_nand4_1 _4667_ (.B(_1095_),
    .C(_1097_),
    .A(_1039_),
    .Y(_1100_),
    .D(_1099_));
 sg13g2_a221oi_1 _4668_ (.B2(net445),
    .C1(_1064_),
    .B1(_0829_),
    .A1(net548),
    .Y(_1101_),
    .A2(_0792_));
 sg13g2_nand2_1 _4669_ (.Y(_1102_),
    .A(_1066_),
    .B(_1101_));
 sg13g2_nor3_1 _4670_ (.A(_2570_),
    .B(_1070_),
    .C(_1071_),
    .Y(_1103_));
 sg13g2_a22oi_1 _4671_ (.Y(_1104_),
    .B1(_0850_),
    .B2(net542),
    .A2(_0842_),
    .A1(_0748_));
 sg13g2_a22oi_1 _4672_ (.Y(_1105_),
    .B1(_2629_),
    .B2(_2639_),
    .A2(net538),
    .A1(_0351_));
 sg13g2_nand4_1 _4673_ (.B(_1103_),
    .C(_1104_),
    .A(_0665_),
    .Y(_1106_),
    .D(_1105_));
 sg13g2_nor4_1 _4674_ (.A(_0318_),
    .B(_0696_),
    .C(_0706_),
    .D(_0795_),
    .Y(_1107_));
 sg13g2_a21oi_1 _4675_ (.A1(net523),
    .A2(_0851_),
    .Y(_1108_),
    .B1(_1062_));
 sg13g2_a22oi_1 _4676_ (.Y(_1110_),
    .B1(_1081_),
    .B2(_0764_),
    .A2(_0847_),
    .A1(_0733_));
 sg13g2_nand4_1 _4677_ (.B(_1107_),
    .C(_1108_),
    .A(_1069_),
    .Y(_1111_),
    .D(_1110_));
 sg13g2_nor4_1 _4678_ (.A(_1100_),
    .B(_1102_),
    .C(_1106_),
    .D(_1111_),
    .Y(_1112_));
 sg13g2_and4_1 _4679_ (.A(_1034_),
    .B(_1058_),
    .C(_1093_),
    .D(_1112_),
    .X(_1113_));
 sg13g2_nand4_1 _4680_ (.B(_1091_),
    .C(_1092_),
    .A(_1046_),
    .Y(_1114_),
    .D(_1113_));
 sg13g2_nor4_1 _4681_ (.A(_1050_),
    .B(_1060_),
    .C(_1083_),
    .D(_1114_),
    .Y(_1115_));
 sg13g2_a21oi_1 _4682_ (.A1(_0641_),
    .A2(_1002_),
    .Y(_1116_),
    .B1(_0299_));
 sg13g2_o21ai_1 _4683_ (.B1(_0255_),
    .Y(_1117_),
    .A1(_0575_),
    .A2(_1116_));
 sg13g2_nor2b_1 _4684_ (.A(_0620_),
    .B_N(_1117_),
    .Y(_1118_));
 sg13g2_nand2_1 _4685_ (.Y(_1119_),
    .A(_0681_),
    .B(_0566_));
 sg13g2_nand2_1 _4686_ (.Y(_1121_),
    .A(_0500_),
    .B(_1119_));
 sg13g2_a21oi_1 _4687_ (.A1(net534),
    .A2(_0566_),
    .Y(_1122_),
    .B1(_1121_));
 sg13g2_and2_1 _4688_ (.A(_0587_),
    .B(_1053_),
    .X(_1123_));
 sg13g2_nor3_2 _4689_ (.A(_0164_),
    .B(_0175_),
    .C(net495),
    .Y(_1124_));
 sg13g2_a21oi_1 _4690_ (.A1(_0570_),
    .A2(_0585_),
    .Y(_1125_),
    .B1(_0575_));
 sg13g2_nand2_1 _4691_ (.Y(_1126_),
    .A(_1124_),
    .B(_1125_));
 sg13g2_or2_1 _4692_ (.X(_1127_),
    .B(_1123_),
    .A(_1122_));
 sg13g2_nand2_1 _4693_ (.Y(_1128_),
    .A(_1115_),
    .B(_1126_));
 sg13g2_nor4_1 _4694_ (.A(_1033_),
    .B(_1118_),
    .C(_1127_),
    .D(_1128_),
    .Y(_1129_));
 sg13g2_o21ai_1 _4695_ (.B1(_1129_),
    .Y(_1130_),
    .A1(_0328_),
    .A2(_0421_));
 sg13g2_nor2_1 _4696_ (.A(_0992_),
    .B(_1130_),
    .Y(_1132_));
 sg13g2_a21oi_1 _4697_ (.A1(_1001_),
    .A2(_1132_),
    .Y(uo_out[0]),
    .B1(_0637_));
 sg13g2_nand2_1 _4698_ (.Y(_1133_),
    .A(_0951_),
    .B(_0957_));
 sg13g2_nor4_1 _4699_ (.A(_2448_),
    .B(_0959_),
    .C(_0980_),
    .D(_1133_),
    .Y(_1134_));
 sg13g2_nand2_1 _4700_ (.Y(_1135_),
    .A(net547),
    .B(_0234_));
 sg13g2_nand4_1 _4701_ (.B(net547),
    .C(_1755_),
    .A(_0714_),
    .Y(_1136_),
    .D(_0234_));
 sg13g2_a21oi_1 _4702_ (.A1(net568),
    .A2(_0549_),
    .Y(_1137_),
    .B1(_2587_));
 sg13g2_a21oi_1 _4703_ (.A1(_2031_),
    .A2(_0981_),
    .Y(_1138_),
    .B1(_1134_));
 sg13g2_and4_1 _4704_ (.A(_2639_),
    .B(_1136_),
    .C(_1137_),
    .D(_1138_),
    .X(_1139_));
 sg13g2_xnor2_1 _4705_ (.Y(_1140_),
    .A(net632),
    .B(_2670_));
 sg13g2_a22oi_1 _4706_ (.Y(_1142_),
    .B1(_2669_),
    .B2(net557),
    .A2(_2638_),
    .A1(_2636_));
 sg13g2_nand3b_1 _4707_ (.B(_2638_),
    .C(_1140_),
    .Y(_1143_),
    .A_N(net518));
 sg13g2_o21ai_1 _4708_ (.B1(net518),
    .Y(_1144_),
    .A1(net557),
    .A2(_2669_));
 sg13g2_and2_1 _4709_ (.A(_1143_),
    .B(_1144_),
    .X(_1145_));
 sg13g2_nand3b_1 _4710_ (.B(_2672_),
    .C(_2638_),
    .Y(_1146_),
    .A_N(net518));
 sg13g2_o21ai_1 _4711_ (.B1(_2674_),
    .Y(_1147_),
    .A1(_2639_),
    .A2(net518));
 sg13g2_and2_1 _4712_ (.A(_1146_),
    .B(_1147_),
    .X(_1148_));
 sg13g2_inv_2 _4713_ (.Y(_1149_),
    .A(_1148_));
 sg13g2_nand2_1 _4714_ (.Y(_1150_),
    .A(_1145_),
    .B(_1148_));
 sg13g2_nor2_1 _4715_ (.A(_2036_),
    .B(_0570_),
    .Y(_1151_));
 sg13g2_o21ai_1 _4716_ (.B1(net521),
    .Y(_1153_),
    .A1(net529),
    .A2(_0570_));
 sg13g2_a221oi_1 _4717_ (.B2(net541),
    .C1(_0950_),
    .B1(_0654_),
    .A1(net528),
    .Y(_1154_),
    .A2(_0569_));
 sg13g2_nand3_1 _4718_ (.B(net529),
    .C(net521),
    .A(net596),
    .Y(_1155_));
 sg13g2_o21ai_1 _4719_ (.B1(_1155_),
    .Y(_1156_),
    .A1(_1151_),
    .A2(_1154_));
 sg13g2_and2_1 _4720_ (.A(_1251_),
    .B(_1156_),
    .X(_1157_));
 sg13g2_nand2_2 _4721_ (.Y(_1158_),
    .A(_1251_),
    .B(_1156_));
 sg13g2_o21ai_1 _4722_ (.B1(_2591_),
    .Y(_1159_),
    .A1(net561),
    .A2(_1240_));
 sg13g2_mux2_1 _4723_ (.A0(_2019_),
    .A1(_1159_),
    .S(_0569_),
    .X(_1160_));
 sg13g2_nand2_1 _4724_ (.Y(_1161_),
    .A(_1251_),
    .B(_0583_));
 sg13g2_xnor2_1 _4725_ (.Y(_1162_),
    .A(net582),
    .B(_1161_));
 sg13g2_a21oi_1 _4726_ (.A1(_2572_),
    .A2(_0583_),
    .Y(_1164_),
    .B1(net519));
 sg13g2_a21oi_1 _4727_ (.A1(net519),
    .A2(_1162_),
    .Y(_1165_),
    .B1(_1164_));
 sg13g2_mux2_1 _4728_ (.A0(_0971_),
    .A1(_0969_),
    .S(_1160_),
    .X(_1166_));
 sg13g2_o21ai_1 _4729_ (.B1(_1166_),
    .Y(_1167_),
    .A1(net528),
    .A2(_1165_));
 sg13g2_or2_1 _4730_ (.X(_1168_),
    .B(_1167_),
    .A(_1158_));
 sg13g2_nand4_1 _4731_ (.B(net572),
    .C(net560),
    .A(net562),
    .Y(_1169_),
    .D(_2572_));
 sg13g2_o21ai_1 _4732_ (.B1(_2047_),
    .Y(_1170_),
    .A1(net528),
    .A2(net519));
 sg13g2_and2_1 _4733_ (.A(_0569_),
    .B(_1169_),
    .X(_1171_));
 sg13g2_and2_1 _4734_ (.A(_1170_),
    .B(_1171_),
    .X(_1172_));
 sg13g2_a22oi_1 _4735_ (.Y(_1173_),
    .B1(_1170_),
    .B2(_1171_),
    .A2(_0952_),
    .A1(net532));
 sg13g2_a21o_2 _4736_ (.A2(_0952_),
    .A1(net532),
    .B1(_1172_),
    .X(_1175_));
 sg13g2_a21o_1 _4737_ (.A2(_1161_),
    .A1(_1159_),
    .B1(net521),
    .X(_1176_));
 sg13g2_a21oi_1 _4738_ (.A1(net572),
    .A2(_0621_),
    .Y(_1177_),
    .B1(net528));
 sg13g2_a221oi_1 _4739_ (.B2(_1161_),
    .C1(_0570_),
    .B1(_1159_),
    .A1(net562),
    .Y(_1178_),
    .A2(_2573_));
 sg13g2_a221oi_1 _4740_ (.B2(_1177_),
    .C1(_1178_),
    .B1(_1176_),
    .A1(_0570_),
    .Y(_1179_),
    .A2(_0621_));
 sg13g2_nand2_1 _4741_ (.Y(_1180_),
    .A(_1175_),
    .B(net449));
 sg13g2_nand2_1 _4742_ (.Y(_1181_),
    .A(_1145_),
    .B(_1149_));
 sg13g2_xor2_1 _4743_ (.B(_1180_),
    .A(_1168_),
    .X(_1182_));
 sg13g2_nand2b_1 _4744_ (.Y(_1183_),
    .B(_1182_),
    .A_N(_1181_));
 sg13g2_o21ai_1 _4745_ (.B1(_1183_),
    .Y(_1184_),
    .A1(_1168_),
    .A2(_1180_));
 sg13g2_nor3_1 _4746_ (.A(net632),
    .B(_2639_),
    .C(_2670_),
    .Y(_1186_));
 sg13g2_nor2_1 _4747_ (.A(net518),
    .B(_1186_),
    .Y(_1187_));
 sg13g2_xnor2_1 _4748_ (.Y(_1188_),
    .A(net631),
    .B(_1187_));
 sg13g2_nand2_1 _4749_ (.Y(_1189_),
    .A(_1148_),
    .B(_1188_));
 sg13g2_nor2b_1 _4750_ (.A(_1167_),
    .B_N(_1179_),
    .Y(_1190_));
 sg13g2_xor2_1 _4751_ (.B(net449),
    .A(_1167_),
    .X(_1191_));
 sg13g2_nor2_1 _4752_ (.A(_1175_),
    .B(_1191_),
    .Y(_1192_));
 sg13g2_nand2b_1 _4753_ (.Y(_1193_),
    .B(_1192_),
    .A_N(_1189_));
 sg13g2_xnor2_1 _4754_ (.Y(_1194_),
    .A(_1189_),
    .B(_1192_));
 sg13g2_nand2_1 _4755_ (.Y(_1195_),
    .A(_1184_),
    .B(_1194_));
 sg13g2_xnor2_1 _4756_ (.Y(_1197_),
    .A(_1184_),
    .B(_1194_));
 sg13g2_xor2_1 _4757_ (.B(_1197_),
    .A(_1150_),
    .X(_1198_));
 sg13g2_nor2_1 _4758_ (.A(_1218_),
    .B(_0425_),
    .Y(_1199_));
 sg13g2_mux2_1 _4759_ (.A0(net598),
    .A1(_1199_),
    .S(_1153_),
    .X(_1200_));
 sg13g2_inv_1 _4760_ (.Y(_1201_),
    .A(_1200_));
 sg13g2_nand2_1 _4761_ (.Y(_1202_),
    .A(net449),
    .B(_1200_));
 sg13g2_o21ai_1 _4762_ (.B1(_1202_),
    .Y(_1203_),
    .A1(_1158_),
    .A2(_1175_));
 sg13g2_nor2_1 _4763_ (.A(_2635_),
    .B(_1167_),
    .Y(_1204_));
 sg13g2_nand2_1 _4764_ (.Y(_1205_),
    .A(_1173_),
    .B(_1200_));
 sg13g2_nand2_1 _4765_ (.Y(_1206_),
    .A(_1157_),
    .B(net449));
 sg13g2_nor3_1 _4766_ (.A(_1158_),
    .B(_1175_),
    .C(_1202_),
    .Y(_1208_));
 sg13g2_a21oi_2 _4767_ (.B1(_1208_),
    .Y(_1209_),
    .A2(_1204_),
    .A1(_1203_));
 sg13g2_nor2_1 _4768_ (.A(_1175_),
    .B(_1209_),
    .Y(_1210_));
 sg13g2_o21ai_1 _4769_ (.B1(_1206_),
    .Y(_1211_),
    .A1(_1167_),
    .A2(_1201_));
 sg13g2_nand2_1 _4770_ (.Y(_1212_),
    .A(_1210_),
    .B(_1211_));
 sg13g2_nand3b_1 _4771_ (.B(_2680_),
    .C(_2638_),
    .Y(_1213_),
    .A_N(net518));
 sg13g2_o21ai_1 _4772_ (.B1(_2683_),
    .Y(_1214_),
    .A1(_2639_),
    .A2(net518));
 sg13g2_and2_1 _4773_ (.A(_1213_),
    .B(_1214_),
    .X(_1215_));
 sg13g2_and2_1 _4774_ (.A(net448),
    .B(_1215_),
    .X(_1216_));
 sg13g2_nand2_1 _4775_ (.Y(_1217_),
    .A(net448),
    .B(_1215_));
 sg13g2_nand2_1 _4776_ (.Y(_1219_),
    .A(_1157_),
    .B(_1200_));
 sg13g2_nor2_1 _4777_ (.A(_1168_),
    .B(_1202_),
    .Y(_1220_));
 sg13g2_xnor2_1 _4778_ (.Y(_1221_),
    .A(_1217_),
    .B(_1220_));
 sg13g2_nand3b_1 _4779_ (.B(_2638_),
    .C(_1010_),
    .Y(_1222_),
    .A_N(net518));
 sg13g2_o21ai_1 _4780_ (.B1(net644),
    .Y(_1223_),
    .A1(_2639_),
    .A2(_1142_));
 sg13g2_and2_1 _4781_ (.A(_1222_),
    .B(_1223_),
    .X(_1224_));
 sg13g2_nand2_1 _4782_ (.Y(_1225_),
    .A(_1215_),
    .B(_1224_));
 sg13g2_nand2_1 _4783_ (.Y(_1226_),
    .A(_1145_),
    .B(net448));
 sg13g2_and2_1 _4784_ (.A(_1145_),
    .B(_1224_),
    .X(_1227_));
 sg13g2_nand4_1 _4785_ (.B(_1144_),
    .C(_1222_),
    .A(_1143_),
    .Y(_1228_),
    .D(_1223_));
 sg13g2_a22oi_1 _4786_ (.Y(_1230_),
    .B1(_1224_),
    .B2(net448),
    .A2(_1215_),
    .A1(_1145_));
 sg13g2_a21o_2 _4787_ (.A2(_1227_),
    .A1(_1216_),
    .B1(_1230_),
    .X(_1231_));
 sg13g2_nor2_1 _4788_ (.A(_1149_),
    .B(_1231_),
    .Y(_1232_));
 sg13g2_a21oi_1 _4789_ (.A1(_1216_),
    .A2(_1227_),
    .Y(_1233_),
    .B1(_1232_));
 sg13g2_nor2b_1 _4790_ (.A(_1233_),
    .B_N(_1221_),
    .Y(_1234_));
 sg13g2_xnor2_1 _4791_ (.Y(_1235_),
    .A(_1221_),
    .B(_1233_));
 sg13g2_inv_1 _4792_ (.Y(_1236_),
    .A(_1235_));
 sg13g2_xnor2_1 _4793_ (.Y(_1237_),
    .A(_1210_),
    .B(_1211_));
 sg13g2_o21ai_1 _4794_ (.B1(_1212_),
    .Y(_1238_),
    .A1(_1236_),
    .A2(_1237_));
 sg13g2_xnor2_1 _4795_ (.Y(_1239_),
    .A(_1181_),
    .B(_1182_));
 sg13g2_a21oi_1 _4796_ (.A1(_1216_),
    .A2(_1220_),
    .Y(_1241_),
    .B1(_1234_));
 sg13g2_xnor2_1 _4797_ (.Y(_1242_),
    .A(_1238_),
    .B(_1239_));
 sg13g2_nor2_1 _4798_ (.A(_1241_),
    .B(_1242_),
    .Y(_1243_));
 sg13g2_a21oi_1 _4799_ (.A1(_1238_),
    .A2(_1239_),
    .Y(_1244_),
    .B1(_1243_));
 sg13g2_nor2b_1 _4800_ (.A(_1244_),
    .B_N(_1198_),
    .Y(_1245_));
 sg13g2_xnor2_1 _4801_ (.Y(_1246_),
    .A(_1198_),
    .B(_1244_));
 sg13g2_xnor2_1 _4802_ (.Y(_1247_),
    .A(_1175_),
    .B(_1209_));
 sg13g2_o21ai_1 _4803_ (.B1(_1203_),
    .Y(_1248_),
    .A1(_1205_),
    .A2(_1206_));
 sg13g2_xnor2_1 _4804_ (.Y(_1249_),
    .A(_1204_),
    .B(_1248_));
 sg13g2_nand2b_1 _4805_ (.Y(_1250_),
    .B(_1249_),
    .A_N(_1247_));
 sg13g2_xor2_1 _4806_ (.B(_1249_),
    .A(_1247_),
    .X(_1252_));
 sg13g2_and2_1 _4807_ (.A(_1148_),
    .B(_1215_),
    .X(_1253_));
 sg13g2_nand4_1 _4808_ (.B(_1147_),
    .C(_1213_),
    .A(_1146_),
    .Y(_1254_),
    .D(_1214_));
 sg13g2_nand2_2 _4809_ (.Y(_1255_),
    .A(net647),
    .B(net448));
 sg13g2_xor2_1 _4810_ (.B(_1254_),
    .A(_1228_),
    .X(_1256_));
 sg13g2_nor2b_1 _4811_ (.A(_1255_),
    .B_N(_1256_),
    .Y(_1257_));
 sg13g2_a21oi_2 _4812_ (.B1(_1257_),
    .Y(_1258_),
    .A2(_1253_),
    .A1(_1227_));
 sg13g2_xnor2_1 _4813_ (.Y(_1259_),
    .A(_1148_),
    .B(_1231_));
 sg13g2_nand2b_1 _4814_ (.Y(_1260_),
    .B(_1259_),
    .A_N(_1209_));
 sg13g2_xnor2_1 _4815_ (.Y(_1261_),
    .A(_1209_),
    .B(_1259_));
 sg13g2_inv_1 _4816_ (.Y(_1263_),
    .A(_1261_));
 sg13g2_xor2_1 _4817_ (.B(_1261_),
    .A(_1258_),
    .X(_1264_));
 sg13g2_o21ai_1 _4818_ (.B1(_1250_),
    .Y(_1265_),
    .A1(_1252_),
    .A2(_1264_));
 sg13g2_xor2_1 _4819_ (.B(_1237_),
    .A(_1235_),
    .X(_1266_));
 sg13g2_inv_1 _4820_ (.Y(_1267_),
    .A(_1266_));
 sg13g2_xor2_1 _4821_ (.B(_1266_),
    .A(_1265_),
    .X(_1268_));
 sg13g2_o21ai_1 _4822_ (.B1(_1260_),
    .Y(_1269_),
    .A1(_1258_),
    .A2(_1263_));
 sg13g2_nor2_1 _4823_ (.A(_1217_),
    .B(_1227_),
    .Y(_1270_));
 sg13g2_xnor2_1 _4824_ (.Y(_1271_),
    .A(_1269_),
    .B(_1270_));
 sg13g2_nor2_1 _4825_ (.A(_1268_),
    .B(_1271_),
    .Y(_1272_));
 sg13g2_a21oi_1 _4826_ (.A1(_1265_),
    .A2(_1267_),
    .Y(_1274_),
    .B1(_1272_));
 sg13g2_xor2_1 _4827_ (.B(_1242_),
    .A(_1241_),
    .X(_1275_));
 sg13g2_nor2b_1 _4828_ (.A(_1274_),
    .B_N(_1275_),
    .Y(_1276_));
 sg13g2_xnor2_1 _4829_ (.Y(_1277_),
    .A(_1274_),
    .B(_1275_));
 sg13g2_nor2_1 _4830_ (.A(_1227_),
    .B(_1269_),
    .Y(_1278_));
 sg13g2_nor2_1 _4831_ (.A(_1217_),
    .B(_1278_),
    .Y(_1279_));
 sg13g2_a21oi_1 _4832_ (.A1(_1277_),
    .A2(_1279_),
    .Y(_1280_),
    .B1(_1276_));
 sg13g2_nor2b_1 _4833_ (.A(_1280_),
    .B_N(_1246_),
    .Y(_1281_));
 sg13g2_inv_1 _4834_ (.Y(_1282_),
    .A(_1281_));
 sg13g2_nand2_2 _4835_ (.Y(_1283_),
    .A(net647),
    .B(_1148_));
 sg13g2_nand2_2 _4836_ (.Y(_1285_),
    .A(net647),
    .B(_1145_));
 sg13g2_nand2_1 _4837_ (.Y(_1286_),
    .A(_1148_),
    .B(_1224_));
 sg13g2_nor2_1 _4838_ (.A(_1228_),
    .B(_1283_),
    .Y(_1287_));
 sg13g2_xnor2_1 _4839_ (.Y(_1288_),
    .A(_1255_),
    .B(_1256_));
 sg13g2_xor2_1 _4840_ (.B(_1256_),
    .A(_1255_),
    .X(_1289_));
 sg13g2_nand2_1 _4841_ (.Y(_1290_),
    .A(net602),
    .B(_1173_));
 sg13g2_nand4_1 _4842_ (.B(_1173_),
    .C(net449),
    .A(net602),
    .Y(_1291_),
    .D(_1200_));
 sg13g2_a22oi_1 _4843_ (.Y(_1292_),
    .B1(_1200_),
    .B2(_1173_),
    .A2(net449),
    .A1(net602));
 sg13g2_a21oi_1 _4844_ (.A1(_1158_),
    .A2(_1291_),
    .Y(_1293_),
    .B1(_1292_));
 sg13g2_xnor2_1 _4845_ (.Y(_1294_),
    .A(_1288_),
    .B(_1293_));
 sg13g2_nor3_1 _4846_ (.A(_1228_),
    .B(_1283_),
    .C(_1294_),
    .Y(_1296_));
 sg13g2_xor2_1 _4847_ (.B(_1294_),
    .A(_1287_),
    .X(_1297_));
 sg13g2_o21ai_1 _4848_ (.B1(_1291_),
    .Y(_1298_),
    .A1(_1157_),
    .A2(_1292_));
 sg13g2_nand2b_1 _4849_ (.Y(_1299_),
    .B(_1298_),
    .A_N(_1297_));
 sg13g2_xnor2_1 _4850_ (.Y(_1300_),
    .A(_1252_),
    .B(_1264_));
 sg13g2_nor2_1 _4851_ (.A(_1299_),
    .B(_1300_),
    .Y(_1301_));
 sg13g2_xor2_1 _4852_ (.B(_1300_),
    .A(_1299_),
    .X(_1302_));
 sg13g2_a21o_1 _4853_ (.A2(_1293_),
    .A1(_1288_),
    .B1(_1296_),
    .X(_1303_));
 sg13g2_nand2b_1 _4854_ (.Y(_1304_),
    .B(_1303_),
    .A_N(_1231_));
 sg13g2_xor2_1 _4855_ (.B(_1303_),
    .A(_1231_),
    .X(_1305_));
 sg13g2_xor2_1 _4856_ (.B(_1305_),
    .A(_1258_),
    .X(_1307_));
 sg13g2_a21oi_1 _4857_ (.A1(_1302_),
    .A2(_1307_),
    .Y(_1308_),
    .B1(_1301_));
 sg13g2_xnor2_1 _4858_ (.Y(_1309_),
    .A(_1268_),
    .B(_1271_));
 sg13g2_nor2_1 _4859_ (.A(_1308_),
    .B(_1309_),
    .Y(_1310_));
 sg13g2_o21ai_1 _4860_ (.B1(_1304_),
    .Y(_1311_),
    .A1(_1258_),
    .A2(_1305_));
 sg13g2_xor2_1 _4861_ (.B(_1309_),
    .A(_1308_),
    .X(_1312_));
 sg13g2_a21oi_1 _4862_ (.A1(_1311_),
    .A2(_1312_),
    .Y(_1313_),
    .B1(_1310_));
 sg13g2_xor2_1 _4863_ (.B(_1279_),
    .A(_1277_),
    .X(_1314_));
 sg13g2_nand2b_1 _4864_ (.Y(_1315_),
    .B(_1314_),
    .A_N(_1313_));
 sg13g2_xnor2_1 _4865_ (.Y(_1316_),
    .A(_1157_),
    .B(_1290_));
 sg13g2_xor2_1 _4866_ (.B(_1286_),
    .A(_1285_),
    .X(_1318_));
 sg13g2_nor2b_1 _4867_ (.A(_1219_),
    .B_N(_1318_),
    .Y(_1319_));
 sg13g2_xnor2_1 _4868_ (.Y(_1320_),
    .A(_1219_),
    .B(_1318_));
 sg13g2_nand2_1 _4869_ (.Y(_1321_),
    .A(_1316_),
    .B(_1320_));
 sg13g2_o21ai_1 _4870_ (.B1(_1321_),
    .Y(_1322_),
    .A1(_1158_),
    .A2(_1290_));
 sg13g2_xnor2_1 _4871_ (.Y(_1323_),
    .A(_1297_),
    .B(_1298_));
 sg13g2_nand2_1 _4872_ (.Y(_1324_),
    .A(_1322_),
    .B(_1323_));
 sg13g2_xnor2_1 _4873_ (.Y(_1325_),
    .A(_1322_),
    .B(_1323_));
 sg13g2_xnor2_1 _4874_ (.Y(_1326_),
    .A(_1215_),
    .B(_1286_));
 sg13g2_nand2b_1 _4875_ (.Y(_1327_),
    .B(_1326_),
    .A_N(_1285_));
 sg13g2_o21ai_1 _4876_ (.B1(_1327_),
    .Y(_1329_),
    .A1(_1149_),
    .A2(_1225_));
 sg13g2_xnor2_1 _4877_ (.Y(_1330_),
    .A(_1289_),
    .B(_1319_));
 sg13g2_and2_1 _4878_ (.A(_1329_),
    .B(_1330_),
    .X(_1331_));
 sg13g2_xnor2_1 _4879_ (.Y(_1332_),
    .A(_1329_),
    .B(_1330_));
 sg13g2_o21ai_1 _4880_ (.B1(_1324_),
    .Y(_1333_),
    .A1(_1325_),
    .A2(_1332_));
 sg13g2_xnor2_1 _4881_ (.Y(_1334_),
    .A(_1302_),
    .B(_1307_));
 sg13g2_nor2b_1 _4882_ (.A(_1334_),
    .B_N(_1333_),
    .Y(_1335_));
 sg13g2_a21o_1 _4883_ (.A2(_1319_),
    .A1(_1288_),
    .B1(_1331_),
    .X(_1336_));
 sg13g2_nand2b_1 _4884_ (.Y(_1337_),
    .B(_1334_),
    .A_N(_1333_));
 sg13g2_xor2_1 _4885_ (.B(_1334_),
    .A(_1333_),
    .X(_1338_));
 sg13g2_a21oi_1 _4886_ (.A1(_1336_),
    .A2(_1337_),
    .Y(_1340_),
    .B1(_1335_));
 sg13g2_xnor2_1 _4887_ (.Y(_1341_),
    .A(_1311_),
    .B(_1312_));
 sg13g2_nor2_1 _4888_ (.A(_1340_),
    .B(_1341_),
    .Y(_1342_));
 sg13g2_xnor2_1 _4889_ (.Y(_1343_),
    .A(_1340_),
    .B(_1341_));
 sg13g2_nand2_1 _4890_ (.Y(_1344_),
    .A(net602),
    .B(_1156_));
 sg13g2_or2_1 _4891_ (.X(_1345_),
    .B(_1344_),
    .A(_1283_));
 sg13g2_xnor2_1 _4892_ (.Y(_1346_),
    .A(_1285_),
    .B(_1326_));
 sg13g2_nand2b_1 _4893_ (.Y(_1347_),
    .B(_1346_),
    .A_N(_1345_));
 sg13g2_xnor2_1 _4894_ (.Y(_1348_),
    .A(_1345_),
    .B(_1346_));
 sg13g2_nand2b_1 _4895_ (.Y(_1349_),
    .B(_1348_),
    .A_N(_1225_));
 sg13g2_xnor2_1 _4896_ (.Y(_1351_),
    .A(_1225_),
    .B(_1348_));
 sg13g2_xnor2_1 _4897_ (.Y(_1352_),
    .A(_1316_),
    .B(_1320_));
 sg13g2_inv_1 _4898_ (.Y(_1353_),
    .A(_1352_));
 sg13g2_nand2_1 _4899_ (.Y(_1354_),
    .A(_1351_),
    .B(_1353_));
 sg13g2_xor2_1 _4900_ (.B(_1332_),
    .A(_1325_),
    .X(_1355_));
 sg13g2_nor2b_1 _4901_ (.A(_1354_),
    .B_N(_1355_),
    .Y(_1356_));
 sg13g2_nand2_1 _4902_ (.Y(_1357_),
    .A(_1347_),
    .B(_1349_));
 sg13g2_xnor2_1 _4903_ (.Y(_1358_),
    .A(_1354_),
    .B(_1355_));
 sg13g2_a21o_2 _4904_ (.A2(_1358_),
    .A1(_1357_),
    .B1(_1356_),
    .X(_1359_));
 sg13g2_xnor2_1 _4905_ (.Y(_1360_),
    .A(_1336_),
    .B(_1338_));
 sg13g2_nor2_1 _4906_ (.A(_1359_),
    .B(_1360_),
    .Y(_1362_));
 sg13g2_xnor2_1 _4907_ (.Y(_1363_),
    .A(_1351_),
    .B(_1353_));
 sg13g2_xor2_1 _4908_ (.B(_1344_),
    .A(_1283_),
    .X(_1364_));
 sg13g2_nand3_1 _4909_ (.B(_1200_),
    .C(_1364_),
    .A(net602),
    .Y(_1365_));
 sg13g2_o21ai_1 _4910_ (.B1(net647),
    .Y(_1366_),
    .A1(_1148_),
    .A2(_1215_));
 sg13g2_nand2b_1 _4911_ (.Y(_1367_),
    .B(_1254_),
    .A_N(_1366_));
 sg13g2_a21o_1 _4912_ (.A2(_1200_),
    .A1(net602),
    .B1(_1364_),
    .X(_1368_));
 sg13g2_and2_1 _4913_ (.A(_1365_),
    .B(_1368_),
    .X(_1369_));
 sg13g2_nand2b_1 _4914_ (.Y(_1370_),
    .B(_1369_),
    .A_N(_1367_));
 sg13g2_nand2_1 _4915_ (.Y(_1371_),
    .A(_1365_),
    .B(_1370_));
 sg13g2_nand2b_1 _4916_ (.Y(_1373_),
    .B(_1371_),
    .A_N(_1363_));
 sg13g2_xnor2_1 _4917_ (.Y(_1374_),
    .A(_1363_),
    .B(_1371_));
 sg13g2_a21oi_1 _4918_ (.A1(net647),
    .A2(_1253_),
    .Y(_1375_),
    .B1(_1374_));
 sg13g2_nand3_1 _4919_ (.B(_1253_),
    .C(_1374_),
    .A(net647),
    .Y(_1376_));
 sg13g2_xnor2_1 _4920_ (.Y(_1377_),
    .A(_1367_),
    .B(_1369_));
 sg13g2_nand4_1 _4921_ (.B(_1224_),
    .C(_1376_),
    .A(net651),
    .Y(_1378_),
    .D(_1377_));
 sg13g2_nor2_1 _4922_ (.A(_1375_),
    .B(_1378_),
    .Y(_1379_));
 sg13g2_nand2_1 _4923_ (.Y(_1380_),
    .A(_1373_),
    .B(_1376_));
 sg13g2_xnor2_1 _4924_ (.Y(_1381_),
    .A(_1357_),
    .B(_1358_));
 sg13g2_nor2b_1 _4925_ (.A(_1381_),
    .B_N(_1380_),
    .Y(_1382_));
 sg13g2_xnor2_1 _4926_ (.Y(_1384_),
    .A(_1380_),
    .B(_1381_));
 sg13g2_a221oi_1 _4927_ (.B2(_1384_),
    .C1(_1382_),
    .B1(_1379_),
    .A1(_1359_),
    .Y(_1385_),
    .A2(_1360_));
 sg13g2_xor2_1 _4928_ (.B(_1360_),
    .A(_1359_),
    .X(_1386_));
 sg13g2_nor3_1 _4929_ (.A(_1343_),
    .B(_1362_),
    .C(_1385_),
    .Y(_1387_));
 sg13g2_xnor2_1 _4930_ (.Y(_1388_),
    .A(_1313_),
    .B(_1314_));
 sg13g2_o21ai_1 _4931_ (.B1(_1388_),
    .Y(_1389_),
    .A1(_1342_),
    .A2(_1387_));
 sg13g2_xor2_1 _4932_ (.B(_1280_),
    .A(_1246_),
    .X(_1390_));
 sg13g2_a21o_2 _4933_ (.A2(_1389_),
    .A1(_1315_),
    .B1(_1390_),
    .X(_1391_));
 sg13g2_nand2_1 _4934_ (.Y(_1392_),
    .A(_1173_),
    .B(_1190_));
 sg13g2_nand2_1 _4935_ (.Y(_1393_),
    .A(_1193_),
    .B(_1392_));
 sg13g2_nor2_1 _4936_ (.A(_1167_),
    .B(net449),
    .Y(_1395_));
 sg13g2_nor2b_1 _4937_ (.A(_1145_),
    .B_N(net448),
    .Y(_1396_));
 sg13g2_xnor2_1 _4938_ (.Y(_1397_),
    .A(_1395_),
    .B(_1396_));
 sg13g2_inv_1 _4939_ (.Y(_1398_),
    .A(_1397_));
 sg13g2_xnor2_1 _4940_ (.Y(_1399_),
    .A(_1393_),
    .B(_1398_));
 sg13g2_o21ai_1 _4941_ (.B1(_1195_),
    .Y(_1400_),
    .A1(_1150_),
    .A2(_1197_));
 sg13g2_nor2b_1 _4942_ (.A(_1399_),
    .B_N(_1400_),
    .Y(_1401_));
 sg13g2_xnor2_1 _4943_ (.Y(_1402_),
    .A(_1399_),
    .B(_1400_));
 sg13g2_and2_1 _4944_ (.A(_1245_),
    .B(_1402_),
    .X(_1403_));
 sg13g2_xor2_1 _4945_ (.B(_1402_),
    .A(_1245_),
    .X(_1404_));
 sg13g2_inv_1 _4946_ (.Y(_1406_),
    .A(_1404_));
 sg13g2_a21oi_1 _4947_ (.A1(_1282_),
    .A2(_1391_),
    .Y(_1407_),
    .B1(_1406_));
 sg13g2_nand3_1 _4948_ (.B(_1391_),
    .C(_1406_),
    .A(_1282_),
    .Y(_1408_));
 sg13g2_nor2b_1 _4949_ (.A(_1407_),
    .B_N(_1408_),
    .Y(_1409_));
 sg13g2_nor3_1 _4950_ (.A(_1342_),
    .B(_1387_),
    .C(_1388_),
    .Y(_1410_));
 sg13g2_o21ai_1 _4951_ (.B1(_1343_),
    .Y(_1411_),
    .A1(_1362_),
    .A2(_1385_));
 sg13g2_nor2b_1 _4952_ (.A(_1387_),
    .B_N(_1411_),
    .Y(_1412_));
 sg13g2_xnor2_1 _4953_ (.Y(_1413_),
    .A(_1379_),
    .B(_1384_));
 sg13g2_nor2_1 _4954_ (.A(_1382_),
    .B(_1386_),
    .Y(_1414_));
 sg13g2_nor2_1 _4955_ (.A(_1413_),
    .B(_1414_),
    .Y(_1415_));
 sg13g2_o21ai_1 _4956_ (.B1(_1389_),
    .Y(_1417_),
    .A1(_1412_),
    .A2(_1415_));
 sg13g2_nand3_1 _4957_ (.B(_1389_),
    .C(_1390_),
    .A(_1315_),
    .Y(_1418_));
 sg13g2_nand2_1 _4958_ (.Y(_1419_),
    .A(_1391_),
    .B(_1418_));
 sg13g2_o21ai_1 _4959_ (.B1(_1419_),
    .Y(_1420_),
    .A1(_1410_),
    .A2(_1417_));
 sg13g2_nand3_1 _4960_ (.B(net448),
    .C(_1190_),
    .A(_1145_),
    .Y(_1421_));
 sg13g2_o21ai_1 _4961_ (.B1(_1421_),
    .Y(_1422_),
    .A1(net449),
    .A2(net448));
 sg13g2_a21oi_1 _4962_ (.A1(_1167_),
    .A2(_1226_),
    .Y(_1423_),
    .B1(_1422_));
 sg13g2_a21oi_1 _4963_ (.A1(_1393_),
    .A2(_1398_),
    .Y(_1424_),
    .B1(_1401_));
 sg13g2_inv_1 _4964_ (.Y(_1425_),
    .A(_1424_));
 sg13g2_nand2_1 _4965_ (.Y(_1426_),
    .A(_1423_),
    .B(_1425_));
 sg13g2_xnor2_1 _4966_ (.Y(_1428_),
    .A(_1423_),
    .B(_1424_));
 sg13g2_or3_1 _4967_ (.A(_1403_),
    .B(_1407_),
    .C(_1428_),
    .X(_1429_));
 sg13g2_o21ai_1 _4968_ (.B1(_1429_),
    .Y(_1430_),
    .A1(_1409_),
    .A2(_1420_));
 sg13g2_o21ai_1 _4969_ (.B1(_1428_),
    .Y(_1431_),
    .A1(_1403_),
    .A2(_1407_));
 sg13g2_and3_1 _4970_ (.X(_1432_),
    .A(_1421_),
    .B(_1426_),
    .C(_1431_));
 sg13g2_a21oi_2 _4971_ (.B1(_1139_),
    .Y(_1433_),
    .A2(_1432_),
    .A1(_1430_));
 sg13g2_nand3_1 _4972_ (.B(_0281_),
    .C(_0962_),
    .A(_0277_),
    .Y(_1434_));
 sg13g2_a22oi_1 _4973_ (.Y(_1435_),
    .B1(_0954_),
    .B2(_0955_),
    .A2(_0953_),
    .A1(_0221_));
 sg13g2_o21ai_1 _4974_ (.B1(_1434_),
    .Y(_1436_),
    .A1(_0965_),
    .A2(_1435_));
 sg13g2_nand2_1 _4975_ (.Y(_1437_),
    .A(net641),
    .B(_1427_));
 sg13g2_xnor2_1 _4976_ (.Y(_1439_),
    .A(_2701_),
    .B(_2667_));
 sg13g2_nor2_1 _4977_ (.A(_0964_),
    .B(_1439_),
    .Y(_1440_));
 sg13g2_o21ai_1 _4978_ (.B1(_1436_),
    .Y(_1441_),
    .A1(_0221_),
    .A2(_0953_));
 sg13g2_nand2_1 _4979_ (.Y(_1442_),
    .A(_2556_),
    .B(_2667_));
 sg13g2_nand2b_1 _4980_ (.Y(_1443_),
    .B(_1437_),
    .A_N(net627));
 sg13g2_nand2_1 _4981_ (.Y(_1444_),
    .A(_1442_),
    .B(_1443_));
 sg13g2_a22oi_1 _4982_ (.Y(_1445_),
    .B1(_1444_),
    .B2(_0972_),
    .A2(_1439_),
    .A1(_0964_));
 sg13g2_o21ai_1 _4983_ (.B1(_1445_),
    .Y(_1446_),
    .A1(_1440_),
    .A2(_1441_));
 sg13g2_nand2_1 _4984_ (.Y(_1447_),
    .A(_0234_),
    .B(_1437_));
 sg13g2_xnor2_1 _4985_ (.Y(_1448_),
    .A(net556),
    .B(_1443_));
 sg13g2_o21ai_1 _4986_ (.B1(_1446_),
    .Y(_1450_),
    .A1(_0972_),
    .A2(_1444_));
 sg13g2_a21oi_1 _4987_ (.A1(_0975_),
    .A2(_1448_),
    .Y(_1451_),
    .B1(_1450_));
 sg13g2_nand2_1 _4988_ (.Y(_1452_),
    .A(net619),
    .B(_1447_));
 sg13g2_xnor2_1 _4989_ (.Y(_1453_),
    .A(net554),
    .B(_1447_));
 sg13g2_nand2_1 _4990_ (.Y(_1454_),
    .A(_0244_),
    .B(_1453_));
 sg13g2_o21ai_1 _4991_ (.B1(_1454_),
    .Y(_1455_),
    .A1(_0975_),
    .A2(_1448_));
 sg13g2_nor2_1 _4992_ (.A(_0244_),
    .B(_1453_),
    .Y(_1456_));
 sg13g2_xnor2_1 _4993_ (.Y(_1457_),
    .A(net552),
    .B(_1452_));
 sg13g2_a21oi_1 _4994_ (.A1(_0980_),
    .A2(_1457_),
    .Y(_1458_),
    .B1(_1456_));
 sg13g2_o21ai_1 _4995_ (.B1(_1458_),
    .Y(_1459_),
    .A1(_1451_),
    .A2(_1455_));
 sg13g2_nand2b_1 _4996_ (.Y(_1461_),
    .B(_0982_),
    .A_N(_1452_));
 sg13g2_nand2_1 _4997_ (.Y(_1462_),
    .A(net551),
    .B(_1137_));
 sg13g2_a221oi_1 _4998_ (.B2(_0553_),
    .C1(_1462_),
    .B1(_1442_),
    .A1(net614),
    .Y(_1463_),
    .A2(_0981_));
 sg13g2_nand2_1 _4999_ (.Y(_1464_),
    .A(_2031_),
    .B(_1134_));
 sg13g2_nand4_1 _5000_ (.B(_1461_),
    .C(_1463_),
    .A(_1459_),
    .Y(_1465_),
    .D(_1464_));
 sg13g2_o21ai_1 _5001_ (.B1(_0990_),
    .Y(_1466_),
    .A1(_1433_),
    .A2(_1465_));
 sg13g2_nor2_1 _5002_ (.A(_2573_),
    .B(_0642_),
    .Y(_1467_));
 sg13g2_nand2b_1 _5003_ (.Y(_1468_),
    .B(_1467_),
    .A_N(_0325_));
 sg13g2_a21oi_1 _5004_ (.A1(_1030_),
    .A2(_1468_),
    .Y(_1469_),
    .B1(_0269_));
 sg13g2_nand2b_1 _5005_ (.Y(_1470_),
    .B(_0420_),
    .A_N(_0418_));
 sg13g2_nor2_1 _5006_ (.A(_0410_),
    .B(_0411_),
    .Y(_1472_));
 sg13g2_and2_1 _5007_ (.A(_0414_),
    .B(_1472_),
    .X(_1473_));
 sg13g2_nor4_1 _5008_ (.A(_0404_),
    .B(_0416_),
    .C(_1470_),
    .D(_1473_),
    .Y(_1474_));
 sg13g2_a21o_1 _5009_ (.A2(_1472_),
    .A1(_0416_),
    .B1(_1470_),
    .X(_1475_));
 sg13g2_a22oi_1 _5010_ (.Y(_1476_),
    .B1(_1475_),
    .B2(_0409_),
    .A2(_1474_),
    .A1(_0408_));
 sg13g2_o21ai_1 _5011_ (.B1(net521),
    .Y(_1477_),
    .A1(_0493_),
    .A2(_0658_));
 sg13g2_o21ai_1 _5012_ (.B1(_0576_),
    .Y(_1478_),
    .A1(_0299_),
    .A2(_1467_));
 sg13g2_xnor2_1 _5013_ (.Y(_1479_),
    .A(net622),
    .B(_0956_));
 sg13g2_nor2_1 _5014_ (.A(net475),
    .B(_1479_),
    .Y(_1480_));
 sg13g2_xnor2_1 _5015_ (.Y(_1481_),
    .A(net628),
    .B(net547));
 sg13g2_a22oi_1 _5016_ (.Y(_1483_),
    .B1(net476),
    .B2(_1438_),
    .A2(_2329_),
    .A1(net637));
 sg13g2_o21ai_1 _5017_ (.B1(_1483_),
    .Y(_1484_),
    .A1(_0305_),
    .A2(_0622_));
 sg13g2_or2_1 _5018_ (.X(_1485_),
    .B(_0224_),
    .A(_1438_));
 sg13g2_nor2_1 _5019_ (.A(net586),
    .B(_1481_),
    .Y(_1486_));
 sg13g2_a22oi_1 _5020_ (.Y(_1487_),
    .B1(_1484_),
    .B2(_1485_),
    .A2(_1481_),
    .A1(net586));
 sg13g2_nor3_1 _5021_ (.A(_1480_),
    .B(_1486_),
    .C(_1487_),
    .Y(_1488_));
 sg13g2_xnor2_1 _5022_ (.Y(_1489_),
    .A(net616),
    .B(_1135_));
 sg13g2_a221oi_1 _5023_ (.B2(_0245_),
    .C1(_1488_),
    .B1(_1489_),
    .A1(net475),
    .Y(_1490_),
    .A2(_1479_));
 sg13g2_nor2b_1 _5024_ (.A(_0250_),
    .B_N(_1135_),
    .Y(_1491_));
 sg13g2_or3_1 _5025_ (.A(_0253_),
    .B(_1490_),
    .C(_1491_),
    .X(_1492_));
 sg13g2_a21oi_1 _5026_ (.A1(_1478_),
    .A2(_1492_),
    .Y(_1494_),
    .B1(_0620_));
 sg13g2_and3_1 _5027_ (.X(_1495_),
    .A(_0569_),
    .B(_0576_),
    .C(_1124_));
 sg13g2_nor2_1 _5028_ (.A(net467),
    .B(_0864_),
    .Y(_1496_));
 sg13g2_inv_1 _5029_ (.Y(_1497_),
    .A(_1496_));
 sg13g2_a21oi_1 _5030_ (.A1(net480),
    .A2(net446),
    .Y(_1498_),
    .B1(_1497_));
 sg13g2_o21ai_1 _5031_ (.B1(_0706_),
    .Y(_1499_),
    .A1(_0771_),
    .A2(_1498_));
 sg13g2_nand4_1 _5032_ (.B(_0717_),
    .C(_0770_),
    .A(_0676_),
    .Y(_1500_),
    .D(_0881_));
 sg13g2_a21o_1 _5033_ (.A2(_0891_),
    .A1(_2636_),
    .B1(_2582_),
    .X(_1501_));
 sg13g2_nand3_1 _5034_ (.B(_2584_),
    .C(_1501_),
    .A(_0604_),
    .Y(_1502_));
 sg13g2_a21oi_1 _5035_ (.A1(net629),
    .A2(_0888_),
    .Y(_1503_),
    .B1(_2555_));
 sg13g2_a221oi_1 _5036_ (.B2(net629),
    .C1(_2555_),
    .B1(_0888_),
    .A1(net618),
    .Y(_1505_),
    .A2(_2582_));
 sg13g2_inv_1 _5037_ (.Y(_1506_),
    .A(_1505_));
 sg13g2_a21o_1 _5038_ (.A2(_1506_),
    .A1(_1502_),
    .B1(net606),
    .X(_1507_));
 sg13g2_nand2_1 _5039_ (.Y(_1508_),
    .A(net554),
    .B(_1503_));
 sg13g2_nand4_1 _5040_ (.B(net486),
    .C(_1502_),
    .A(net606),
    .Y(_1509_),
    .D(_1508_));
 sg13g2_nand3_1 _5041_ (.B(_1507_),
    .C(_1509_),
    .A(net456),
    .Y(_1510_));
 sg13g2_a21oi_1 _5042_ (.A1(_0719_),
    .A2(_1510_),
    .Y(_1511_),
    .B1(_0886_));
 sg13g2_nor2_1 _5043_ (.A(_0768_),
    .B(_0865_),
    .Y(_1512_));
 sg13g2_nor2b_1 _5044_ (.A(_1512_),
    .B_N(_0903_),
    .Y(_1513_));
 sg13g2_nor4_1 _5045_ (.A(net619),
    .B(net552),
    .C(net609),
    .D(net525),
    .Y(_1514_));
 sg13g2_o21ai_1 _5046_ (.B1(_0333_),
    .Y(_1516_),
    .A1(net633),
    .A2(_2667_));
 sg13g2_nor2b_1 _5047_ (.A(_1207_),
    .B_N(_2019_),
    .Y(_1517_));
 sg13g2_a221oi_1 _5048_ (.B2(_0747_),
    .C1(net556),
    .B1(_0359_),
    .A1(net627),
    .Y(_1518_),
    .A2(net547));
 sg13g2_o21ai_1 _5049_ (.B1(_1514_),
    .Y(_1519_),
    .A1(_1427_),
    .A2(_0235_));
 sg13g2_o21ai_1 _5050_ (.B1(_1516_),
    .Y(_1520_),
    .A1(net468),
    .A2(_1517_));
 sg13g2_nor4_1 _5051_ (.A(_0569_),
    .B(_1518_),
    .C(_1519_),
    .D(_1520_),
    .Y(_1521_));
 sg13g2_nor3_1 _5052_ (.A(_2553_),
    .B(_2557_),
    .C(_0887_),
    .Y(_1522_));
 sg13g2_nor3_1 _5053_ (.A(_2447_),
    .B(_2573_),
    .C(_0597_),
    .Y(_1523_));
 sg13g2_nor2_1 _5054_ (.A(_0494_),
    .B(_1523_),
    .Y(_1524_));
 sg13g2_a21oi_1 _5055_ (.A1(_0934_),
    .A2(_2642_),
    .Y(_1525_),
    .B1(_2594_));
 sg13g2_nor2b_1 _5056_ (.A(_0712_),
    .B_N(net577),
    .Y(_1527_));
 sg13g2_nor4_1 _5057_ (.A(net606),
    .B(_1109_),
    .C(_1079_),
    .D(_1525_),
    .Y(_1528_));
 sg13g2_o21ai_1 _5058_ (.B1(_1528_),
    .Y(_1529_),
    .A1(net614),
    .A2(_1522_));
 sg13g2_nor3_1 _5059_ (.A(_1524_),
    .B(_1527_),
    .C(_1529_),
    .Y(_1530_));
 sg13g2_o21ai_1 _5060_ (.B1(_0988_),
    .Y(_1531_),
    .A1(_1521_),
    .A2(_1530_));
 sg13g2_nand2_1 _5061_ (.Y(_1532_),
    .A(net524),
    .B(_0612_));
 sg13g2_nand2_1 _5062_ (.Y(_1533_),
    .A(net527),
    .B(_1532_));
 sg13g2_nand4_1 _5063_ (.B(_0439_),
    .C(_0498_),
    .A(_0131_),
    .Y(_1534_),
    .D(_0617_));
 sg13g2_o21ai_1 _5064_ (.B1(_0772_),
    .Y(_1535_),
    .A1(_0771_),
    .A2(_0865_));
 sg13g2_o21ai_1 _5065_ (.B1(net482),
    .Y(_1536_),
    .A1(_0602_),
    .A2(net452));
 sg13g2_nand3_1 _5066_ (.B(_0944_),
    .C(_1536_),
    .A(_0942_),
    .Y(_1538_));
 sg13g2_o21ai_1 _5067_ (.B1(_0786_),
    .Y(_1539_),
    .A1(_0651_),
    .A2(_0797_));
 sg13g2_a21oi_1 _5068_ (.A1(net537),
    .A2(_0825_),
    .Y(_1540_),
    .B1(net520));
 sg13g2_nor4_1 _5069_ (.A(_0274_),
    .B(net472),
    .C(_1036_),
    .D(_1540_),
    .Y(_1541_));
 sg13g2_a21oi_1 _5070_ (.A1(_2614_),
    .A2(_1539_),
    .Y(_1542_),
    .B1(_1541_));
 sg13g2_o21ai_1 _5071_ (.B1(_0787_),
    .Y(_1543_),
    .A1(net532),
    .A2(net481));
 sg13g2_nand2_1 _5072_ (.Y(_1544_),
    .A(_0860_),
    .B(_1543_));
 sg13g2_nand3_1 _5073_ (.B(net468),
    .C(_1544_),
    .A(net522),
    .Y(_1545_));
 sg13g2_nor2_1 _5074_ (.A(net486),
    .B(net524),
    .Y(_1546_));
 sg13g2_o21ai_1 _5075_ (.B1(_0753_),
    .Y(_1547_),
    .A1(_1533_),
    .A2(_1546_));
 sg13g2_nand2_1 _5076_ (.Y(_1549_),
    .A(net492),
    .B(_0754_));
 sg13g2_nand3_1 _5077_ (.B(_1547_),
    .C(_1549_),
    .A(_0818_),
    .Y(_1550_));
 sg13g2_nor4_1 _5078_ (.A(_0680_),
    .B(_0734_),
    .C(_0792_),
    .D(_1077_),
    .Y(_1551_));
 sg13g2_nand2_1 _5079_ (.Y(_1552_),
    .A(_0693_),
    .B(net444));
 sg13g2_o21ai_1 _5080_ (.B1(_1552_),
    .Y(_1553_),
    .A1(_0748_),
    .A2(_1551_));
 sg13g2_nor2b_1 _5081_ (.A(_2578_),
    .B_N(_2590_),
    .Y(_1554_));
 sg13g2_a21oi_1 _5082_ (.A1(net489),
    .A2(_0658_),
    .Y(_1555_),
    .B1(net534));
 sg13g2_o21ai_1 _5083_ (.B1(_1555_),
    .Y(_1556_),
    .A1(net489),
    .A2(_0658_));
 sg13g2_a21o_1 _5084_ (.A2(net489),
    .A1(net535),
    .B1(_1555_),
    .X(_1557_));
 sg13g2_a22oi_1 _5085_ (.Y(_1558_),
    .B1(_1557_),
    .B2(_0742_),
    .A2(_1556_),
    .A1(_0741_));
 sg13g2_nor2_1 _5086_ (.A(net519),
    .B(_1558_),
    .Y(_1560_));
 sg13g2_a21oi_1 _5087_ (.A1(_0605_),
    .A2(net450),
    .Y(_1561_),
    .B1(net452));
 sg13g2_nand2b_1 _5088_ (.Y(_1562_),
    .B(_0926_),
    .A_N(_1561_));
 sg13g2_nor4_1 _5089_ (.A(_0340_),
    .B(net538),
    .C(_2573_),
    .D(net473),
    .Y(_1563_));
 sg13g2_nand3_1 _5090_ (.B(_0687_),
    .C(_0844_),
    .A(_0614_),
    .Y(_1564_));
 sg13g2_nand3_1 _5091_ (.B(_1273_),
    .C(_0592_),
    .A(_1131_),
    .Y(_1565_));
 sg13g2_nand2_1 _5092_ (.Y(_1566_),
    .A(net545),
    .B(_1565_));
 sg13g2_nand3_1 _5093_ (.B(_0917_),
    .C(_1566_),
    .A(net534),
    .Y(_1567_));
 sg13g2_o21ai_1 _5094_ (.B1(net453),
    .Y(_1568_),
    .A1(net446),
    .A2(_0768_));
 sg13g2_nand3_1 _5095_ (.B(_0875_),
    .C(_1568_),
    .A(_0688_),
    .Y(_1569_));
 sg13g2_nor2_1 _5096_ (.A(net492),
    .B(net523),
    .Y(_1571_));
 sg13g2_nand2_1 _5097_ (.Y(_1572_),
    .A(net483),
    .B(net542));
 sg13g2_nor2_1 _5098_ (.A(net531),
    .B(_0682_),
    .Y(_1573_));
 sg13g2_nand3_1 _5099_ (.B(_0658_),
    .C(_0739_),
    .A(_0655_),
    .Y(_1574_));
 sg13g2_nand4_1 _5100_ (.B(net526),
    .C(_0700_),
    .A(_0351_),
    .Y(_1575_),
    .D(_0806_));
 sg13g2_nor2_1 _5101_ (.A(net526),
    .B(net483),
    .Y(_1576_));
 sg13g2_nand3b_1 _5102_ (.B(_0811_),
    .C(_0855_),
    .Y(_1577_),
    .A_N(_1576_));
 sg13g2_nand2_1 _5103_ (.Y(_1578_),
    .A(_0580_),
    .B(_0795_));
 sg13g2_a21oi_1 _5104_ (.A1(net484),
    .A2(_0660_),
    .Y(_1579_),
    .B1(_0697_));
 sg13g2_nand3_1 _5105_ (.B(_0752_),
    .C(_0850_),
    .A(_2590_),
    .Y(_1580_));
 sg13g2_nand3_1 _5106_ (.B(_2629_),
    .C(_2638_),
    .A(net491),
    .Y(_1582_));
 sg13g2_nand3b_1 _5107_ (.B(_0580_),
    .C(_0829_),
    .Y(_1583_),
    .A_N(_2608_));
 sg13g2_a22oi_1 _5108_ (.Y(_1584_),
    .B1(_0754_),
    .B2(_0351_),
    .A2(_0661_),
    .A1(_0587_));
 sg13g2_nand3_1 _5109_ (.B(net445),
    .C(_0842_),
    .A(net484),
    .Y(_1585_));
 sg13g2_a21oi_1 _5110_ (.A1(_2582_),
    .A2(net523),
    .Y(_1586_),
    .B1(_0751_));
 sg13g2_nor2b_1 _5111_ (.A(_1586_),
    .B_N(_1070_),
    .Y(_1587_));
 sg13g2_nand2_1 _5112_ (.Y(_1588_),
    .A(net492),
    .B(net445));
 sg13g2_nand3_1 _5113_ (.B(_0746_),
    .C(_0800_),
    .A(net492),
    .Y(_1589_));
 sg13g2_a21oi_1 _5114_ (.A1(net450),
    .A2(_0871_),
    .Y(_1590_),
    .B1(_0771_));
 sg13g2_o21ai_1 _5115_ (.B1(_0614_),
    .Y(_1591_),
    .A1(net490),
    .A2(_0605_));
 sg13g2_a21oi_1 _5116_ (.A1(net490),
    .A2(_0716_),
    .Y(_1593_),
    .B1(_1591_));
 sg13g2_nand2_1 _5117_ (.Y(_1594_),
    .A(_0318_),
    .B(net450));
 sg13g2_a21oi_1 _5118_ (.A1(net480),
    .A2(net455),
    .Y(_1595_),
    .B1(_0715_));
 sg13g2_a21oi_1 _5119_ (.A1(_0775_),
    .A2(_1595_),
    .Y(_1596_),
    .B1(_1594_));
 sg13g2_a21oi_1 _5120_ (.A1(net577),
    .A2(_1042_),
    .Y(_1597_),
    .B1(net573));
 sg13g2_or2_1 _5121_ (.X(_1598_),
    .B(_1597_),
    .A(_0914_));
 sg13g2_a21oi_1 _5122_ (.A1(net543),
    .A2(_0913_),
    .Y(_1599_),
    .B1(net530));
 sg13g2_nor2_1 _5123_ (.A(net486),
    .B(_0855_),
    .Y(_1600_));
 sg13g2_a21o_1 _5124_ (.A2(_1599_),
    .A1(_1598_),
    .B1(_0940_),
    .X(_1601_));
 sg13g2_o21ai_1 _5125_ (.B1(_1045_),
    .Y(_1602_),
    .A1(_1600_),
    .A2(_1601_));
 sg13g2_nor2_1 _5126_ (.A(_0909_),
    .B(_1593_),
    .Y(_1604_));
 sg13g2_a21oi_1 _5127_ (.A1(_0274_),
    .A2(net457),
    .Y(_1605_),
    .B1(net469));
 sg13g2_nor3_1 _5128_ (.A(_0867_),
    .B(_0910_),
    .C(_1605_),
    .Y(_1606_));
 sg13g2_o21ai_1 _5129_ (.B1(_1531_),
    .Y(_1607_),
    .A1(_0719_),
    .A2(_1606_));
 sg13g2_a22oi_1 _5130_ (.Y(_1608_),
    .B1(_1062_),
    .B2(net468),
    .A2(_0916_),
    .A1(net526));
 sg13g2_o21ai_1 _5131_ (.B1(_0285_),
    .Y(_1609_),
    .A1(_0751_),
    .A2(net464));
 sg13g2_nand2_1 _5132_ (.Y(_1610_),
    .A(_0739_),
    .B(_1053_));
 sg13g2_a21oi_1 _5133_ (.A1(net543),
    .A2(_0677_),
    .Y(_1611_),
    .B1(_1587_));
 sg13g2_a21oi_1 _5134_ (.A1(net527),
    .A2(_1554_),
    .Y(_1612_),
    .B1(_1579_));
 sg13g2_nand3_1 _5135_ (.B(_0752_),
    .C(_1532_),
    .A(_0749_),
    .Y(_1613_));
 sg13g2_a21oi_1 _5136_ (.A1(net493),
    .A2(net524),
    .Y(_1615_),
    .B1(_1613_));
 sg13g2_a21o_1 _5137_ (.A2(_1533_),
    .A1(_0831_),
    .B1(_1615_),
    .X(_1616_));
 sg13g2_a21oi_1 _5138_ (.A1(_0646_),
    .A2(_1075_),
    .Y(_1617_),
    .B1(_1563_));
 sg13g2_nand3_1 _5139_ (.B(_1564_),
    .C(_1617_),
    .A(_0849_),
    .Y(_1618_));
 sg13g2_mux2_1 _5140_ (.A0(_0789_),
    .A1(_0805_),
    .S(net451),
    .X(_1619_));
 sg13g2_nand3_1 _5141_ (.B(_1580_),
    .C(_1619_),
    .A(_0652_),
    .Y(_1620_));
 sg13g2_nand3_1 _5142_ (.B(_1584_),
    .C(_1589_),
    .A(_1578_),
    .Y(_1621_));
 sg13g2_nor4_1 _5143_ (.A(_0675_),
    .B(_1618_),
    .C(_1620_),
    .D(_1621_),
    .Y(_1622_));
 sg13g2_nand3_1 _5144_ (.B(_1569_),
    .C(_1622_),
    .A(_1534_),
    .Y(_1623_));
 sg13g2_a21oi_2 _5145_ (.B1(_1623_),
    .Y(_1624_),
    .A2(_1616_),
    .A1(_0753_));
 sg13g2_a22oi_1 _5146_ (.Y(_1626_),
    .B1(_1600_),
    .B2(_0921_),
    .A2(_1573_),
    .A1(_1571_));
 sg13g2_a22oi_1 _5147_ (.Y(_1627_),
    .B1(_0828_),
    .B2(_0578_),
    .A2(_0751_),
    .A1(_0384_));
 sg13g2_nand3_1 _5148_ (.B(_1609_),
    .C(_1627_),
    .A(_1574_),
    .Y(_1628_));
 sg13g2_nand3_1 _5149_ (.B(_1577_),
    .C(_1608_),
    .A(_1567_),
    .Y(_1629_));
 sg13g2_nor4_1 _5150_ (.A(_0815_),
    .B(_0905_),
    .C(_1628_),
    .D(_1629_),
    .Y(_1630_));
 sg13g2_nand4_1 _5151_ (.B(_1575_),
    .C(_1626_),
    .A(_0929_),
    .Y(_1631_),
    .D(_1630_));
 sg13g2_nor4_1 _5152_ (.A(_1513_),
    .B(_1596_),
    .C(_1607_),
    .D(_1631_),
    .Y(_1632_));
 sg13g2_o21ai_1 _5153_ (.B1(_1499_),
    .Y(_1633_),
    .A1(_0883_),
    .A2(_1590_));
 sg13g2_o21ai_1 _5154_ (.B1(_1545_),
    .Y(_1634_),
    .A1(_0329_),
    .A2(_0770_));
 sg13g2_nand4_1 _5155_ (.B(_1585_),
    .C(_1611_),
    .A(_1582_),
    .Y(_1635_),
    .D(_1612_));
 sg13g2_nor4_1 _5156_ (.A(_0672_),
    .B(_1553_),
    .C(_1634_),
    .D(_1635_),
    .Y(_1637_));
 sg13g2_nand4_1 _5157_ (.B(_1550_),
    .C(_1583_),
    .A(_0731_),
    .Y(_1638_),
    .D(_1637_));
 sg13g2_nor3_1 _5158_ (.A(_1560_),
    .B(_1633_),
    .C(_1638_),
    .Y(_1639_));
 sg13g2_a22oi_1 _5159_ (.Y(_1640_),
    .B1(_1604_),
    .B2(_0770_),
    .A2(_1049_),
    .A1(_0776_));
 sg13g2_nand3_1 _5160_ (.B(_1535_),
    .C(_1640_),
    .A(_1500_),
    .Y(_1641_));
 sg13g2_nand4_1 _5161_ (.B(_1542_),
    .C(_1562_),
    .A(_1538_),
    .Y(_1642_),
    .D(_1602_));
 sg13g2_nor4_1 _5162_ (.A(_1495_),
    .B(_1511_),
    .C(_1641_),
    .D(_1642_),
    .Y(_1643_));
 sg13g2_nand4_1 _5163_ (.B(_1632_),
    .C(_1639_),
    .A(_1624_),
    .Y(_1644_),
    .D(_1643_));
 sg13g2_nor3_1 _5164_ (.A(_0567_),
    .B(_1494_),
    .C(_1644_),
    .Y(_1645_));
 sg13g2_o21ai_1 _5165_ (.B1(_1645_),
    .Y(_1646_),
    .A1(_0497_),
    .A2(_1477_));
 sg13g2_a221oi_1 _5166_ (.B2(_0330_),
    .C1(_1646_),
    .B1(_1476_),
    .A1(_0262_),
    .Y(_1648_),
    .A2(_1469_));
 sg13g2_o21ai_1 _5167_ (.B1(_1648_),
    .Y(_1649_),
    .A1(_0987_),
    .A2(_1466_));
 sg13g2_nor2_1 _5168_ (.A(_1000_),
    .B(_1649_),
    .Y(_1650_));
 sg13g2_nand3_1 _5169_ (.B(_2544_),
    .C(_2618_),
    .A(_2745_),
    .Y(_1651_));
 sg13g2_a21o_1 _5170_ (.A2(_1651_),
    .A1(_1766_),
    .B1(_2622_),
    .X(_1652_));
 sg13g2_nand2_1 _5171_ (.Y(_1653_),
    .A(net608),
    .B(net491));
 sg13g2_and3_1 _5172_ (.X(_1654_),
    .A(_2629_),
    .B(_2639_),
    .C(_1653_));
 sg13g2_nor2_1 _5173_ (.A(_2569_),
    .B(_2601_),
    .Y(_1655_));
 sg13g2_a221oi_1 _5174_ (.B2(_1654_),
    .C1(_1655_),
    .B1(_1652_),
    .A1(_2571_),
    .Y(_1656_),
    .A2(net491));
 sg13g2_a21oi_1 _5175_ (.A1(_1650_),
    .A2(_1656_),
    .Y(uo_out[5]),
    .B1(_0637_));
 sg13g2_a21o_1 _5176_ (.A2(_2610_),
    .A1(_2600_),
    .B1(_2601_),
    .X(_1658_));
 sg13g2_a221oi_1 _5177_ (.B2(_2618_),
    .C1(net609),
    .B1(_2544_),
    .A1(net555),
    .Y(_1659_),
    .A2(net553));
 sg13g2_o21ai_1 _5178_ (.B1(_1653_),
    .Y(_1660_),
    .A1(net491),
    .A2(_2639_));
 sg13g2_o21ai_1 _5179_ (.B1(_2629_),
    .Y(_1661_),
    .A1(_1659_),
    .A2(_1660_));
 sg13g2_nor2_1 _5180_ (.A(net524),
    .B(_0754_),
    .Y(_1662_));
 sg13g2_nand2_1 _5181_ (.Y(_1663_),
    .A(net542),
    .B(_0753_));
 sg13g2_o21ai_1 _5182_ (.B1(_0641_),
    .Y(_1664_),
    .A1(_0325_),
    .A2(_1663_));
 sg13g2_and3_1 _5183_ (.X(_1665_),
    .A(_0262_),
    .B(_0268_),
    .C(_1664_));
 sg13g2_nor2_1 _5184_ (.A(_0328_),
    .B(_1476_),
    .Y(_1666_));
 sg13g2_a21oi_1 _5185_ (.A1(_0641_),
    .A2(_1662_),
    .Y(_1667_),
    .B1(_0575_));
 sg13g2_nor2_1 _5186_ (.A(_0620_),
    .B(_1667_),
    .Y(_1669_));
 sg13g2_nand3_1 _5187_ (.B(_2565_),
    .C(_1125_),
    .A(_0219_),
    .Y(_1670_));
 sg13g2_nand2_1 _5188_ (.Y(_1671_),
    .A(_2575_),
    .B(_0987_));
 sg13g2_nand2_1 _5189_ (.Y(_1672_),
    .A(_0990_),
    .B(_1671_));
 sg13g2_and2_1 _5190_ (.A(_0706_),
    .B(_0873_),
    .X(_1673_));
 sg13g2_nand3_1 _5191_ (.B(_0881_),
    .C(_1673_),
    .A(net454),
    .Y(_1674_));
 sg13g2_or2_1 _5192_ (.X(_1675_),
    .B(_1597_),
    .A(_0933_));
 sg13g2_nand2_1 _5193_ (.Y(_1676_),
    .A(net525),
    .B(_1675_));
 sg13g2_nand2_1 _5194_ (.Y(_1677_),
    .A(_1045_),
    .B(_1676_));
 sg13g2_a21oi_1 _5195_ (.A1(_0939_),
    .A2(_1598_),
    .Y(_1678_),
    .B1(_1044_));
 sg13g2_nand2b_1 _5196_ (.Y(_1680_),
    .B(_0915_),
    .A_N(_1678_));
 sg13g2_a21oi_1 _5197_ (.A1(_0732_),
    .A2(_1572_),
    .Y(_1681_),
    .B1(_2606_));
 sg13g2_nor3_1 _5198_ (.A(_2608_),
    .B(_0797_),
    .C(_1074_),
    .Y(_1682_));
 sg13g2_a21oi_1 _5199_ (.A1(net485),
    .A2(_0754_),
    .Y(_1683_),
    .B1(_0819_));
 sg13g2_nand2_1 _5200_ (.Y(_1684_),
    .A(_0851_),
    .B(_0855_));
 sg13g2_a21oi_1 _5201_ (.A1(net488),
    .A2(_0716_),
    .Y(_1685_),
    .B1(_0909_));
 sg13g2_nand2_1 _5202_ (.Y(_1686_),
    .A(_2614_),
    .B(_0858_));
 sg13g2_o21ai_1 _5203_ (.B1(net522),
    .Y(_1687_),
    .A1(net549),
    .A2(net493));
 sg13g2_a22oi_1 _5204_ (.Y(_1688_),
    .B1(_0787_),
    .B2(net549),
    .A2(_0667_),
    .A1(net535));
 sg13g2_nor3_1 _5205_ (.A(net523),
    .B(net479),
    .C(_0668_),
    .Y(_1689_));
 sg13g2_a21oi_1 _5206_ (.A1(_0822_),
    .A2(_1566_),
    .Y(_1691_),
    .B1(_0664_));
 sg13g2_nor2_1 _5207_ (.A(_0870_),
    .B(_1040_),
    .Y(_1692_));
 sg13g2_nor2_1 _5208_ (.A(net444),
    .B(_1692_),
    .Y(_1693_));
 sg13g2_and3_1 _5209_ (.X(_1694_),
    .A(net455),
    .B(_0688_),
    .C(_0709_));
 sg13g2_nor3_1 _5210_ (.A(_0461_),
    .B(_0772_),
    .C(_0900_),
    .Y(_1695_));
 sg13g2_nor3_1 _5211_ (.A(_0600_),
    .B(_0771_),
    .C(_1695_),
    .Y(_1696_));
 sg13g2_o21ai_1 _5212_ (.B1(net487),
    .Y(_1697_),
    .A1(_0602_),
    .A2(_0610_));
 sg13g2_nand2_1 _5213_ (.Y(_1698_),
    .A(_0942_),
    .B(_1697_));
 sg13g2_nand2b_1 _5214_ (.Y(_1699_),
    .B(_1072_),
    .A_N(_0928_));
 sg13g2_nand2b_1 _5215_ (.Y(_1700_),
    .B(_1699_),
    .A_N(net444));
 sg13g2_nor4_2 _5216_ (.A(_0164_),
    .B(_0197_),
    .C(net478),
    .Y(_1702_),
    .D(_1055_));
 sg13g2_a21oi_1 _5217_ (.A1(_0799_),
    .A2(_0860_),
    .Y(_1703_),
    .B1(_0560_));
 sg13g2_nand3_1 _5218_ (.B(_0646_),
    .C(_0795_),
    .A(net549),
    .Y(_1704_));
 sg13g2_nand3b_1 _5219_ (.B(_0848_),
    .C(_1704_),
    .Y(_1705_),
    .A_N(_0792_));
 sg13g2_nand3_1 _5220_ (.B(_2614_),
    .C(_0829_),
    .A(net548),
    .Y(_1706_));
 sg13g2_o21ai_1 _5221_ (.B1(_0850_),
    .Y(_1707_),
    .A1(net484),
    .A2(net464));
 sg13g2_o21ai_1 _5222_ (.B1(_1707_),
    .Y(_1708_),
    .A1(_0395_),
    .A2(net464));
 sg13g2_o21ai_1 _5223_ (.B1(_0917_),
    .Y(_1709_),
    .A1(_1036_),
    .A2(_1053_));
 sg13g2_nand3_1 _5224_ (.B(_0770_),
    .C(_0775_),
    .A(_0318_),
    .Y(_1710_));
 sg13g2_a22oi_1 _5225_ (.Y(_1711_),
    .B1(_1070_),
    .B2(_1586_),
    .A2(_0753_),
    .A1(_0351_));
 sg13g2_nor4_1 _5226_ (.A(_1694_),
    .B(_1702_),
    .C(_1703_),
    .D(_1705_),
    .Y(_1713_));
 sg13g2_a22oi_1 _5227_ (.Y(_1714_),
    .B1(_1071_),
    .B2(_0733_),
    .A2(_0855_),
    .A1(_0851_));
 sg13g2_o21ai_1 _5228_ (.B1(_1677_),
    .Y(_1715_),
    .A1(_0694_),
    .A2(_0927_));
 sg13g2_nor3_1 _5229_ (.A(_1685_),
    .B(_1693_),
    .C(_1696_),
    .Y(_1716_));
 sg13g2_o21ai_1 _5230_ (.B1(_1716_),
    .Y(_1717_),
    .A1(net451),
    .A2(_1691_));
 sg13g2_a22oi_1 _5231_ (.Y(_1718_),
    .B1(_0800_),
    .B2(_1681_),
    .A2(_0741_),
    .A1(net538));
 sg13g2_nand3_1 _5232_ (.B(_1714_),
    .C(_1718_),
    .A(_1711_),
    .Y(_1719_));
 sg13g2_a221oi_1 _5233_ (.B2(_0285_),
    .C1(_1719_),
    .B1(_1576_),
    .A1(_0645_),
    .Y(_1720_),
    .A2(_0646_));
 sg13g2_nor3_1 _5234_ (.A(_1682_),
    .B(_1683_),
    .C(_1689_),
    .Y(_1721_));
 sg13g2_a22oi_1 _5235_ (.Y(_1722_),
    .B1(_1662_),
    .B2(_0814_),
    .A2(_0828_),
    .A1(net522));
 sg13g2_a22oi_1 _5236_ (.Y(_1724_),
    .B1(_1687_),
    .B2(_0810_),
    .A2(_1686_),
    .A1(_0781_));
 sg13g2_nand4_1 _5237_ (.B(_1721_),
    .C(_1722_),
    .A(_1720_),
    .Y(_1725_),
    .D(_1724_));
 sg13g2_or3_1 _5238_ (.A(_1715_),
    .B(_1717_),
    .C(_1725_),
    .X(_1726_));
 sg13g2_nand4_1 _5239_ (.B(_1680_),
    .C(_1700_),
    .A(_1674_),
    .Y(_1727_),
    .D(_1710_));
 sg13g2_nor3_1 _5240_ (.A(_0811_),
    .B(_0831_),
    .C(_0910_),
    .Y(_1728_));
 sg13g2_nand4_1 _5241_ (.B(_0789_),
    .C(_1610_),
    .A(_0678_),
    .Y(_1729_),
    .D(_1728_));
 sg13g2_nor4_1 _5242_ (.A(_0680_),
    .B(_0696_),
    .C(_0745_),
    .D(_0842_),
    .Y(_1730_));
 sg13g2_a221oi_1 _5243_ (.B2(net526),
    .C1(_1123_),
    .B1(_0921_),
    .A1(_0749_),
    .Y(_1731_),
    .A2(_0750_));
 sg13g2_nor2b_1 _5244_ (.A(_1573_),
    .B_N(_1731_),
    .Y(_1732_));
 sg13g2_nand3_1 _5245_ (.B(_1730_),
    .C(_1732_),
    .A(_1688_),
    .Y(_1733_));
 sg13g2_a22oi_1 _5246_ (.Y(_1735_),
    .B1(_1082_),
    .B2(_0764_),
    .A2(_0844_),
    .A1(_0708_));
 sg13g2_nand4_1 _5247_ (.B(_1709_),
    .C(_1713_),
    .A(_1706_),
    .Y(_1736_),
    .D(_1735_));
 sg13g2_nor4_1 _5248_ (.A(_1708_),
    .B(_1729_),
    .C(_1733_),
    .D(_1736_),
    .Y(_1737_));
 sg13g2_nand4_1 _5249_ (.B(_1531_),
    .C(_1698_),
    .A(_1058_),
    .Y(_1738_),
    .D(_1737_));
 sg13g2_nor4_1 _5250_ (.A(_0577_),
    .B(_1726_),
    .C(_1727_),
    .D(_1738_),
    .Y(_1739_));
 sg13g2_nand4_1 _5251_ (.B(_1670_),
    .C(_1672_),
    .A(_1121_),
    .Y(_1740_),
    .D(_1739_));
 sg13g2_nor4_1 _5252_ (.A(_1665_),
    .B(_1666_),
    .C(_1669_),
    .D(_1740_),
    .Y(_1741_));
 sg13g2_nand4_1 _5253_ (.B(_1658_),
    .C(_1661_),
    .A(_2593_),
    .Y(_1742_),
    .D(_1741_));
 sg13g2_nor2b_1 _5254_ (.A(_0637_),
    .B_N(_1742_),
    .Y(uo_out[1]));
 sg13g2_or3_1 _5255_ (.A(net608),
    .B(_2594_),
    .C(_2622_),
    .X(_1743_));
 sg13g2_nand3_1 _5256_ (.B(_1654_),
    .C(_1743_),
    .A(_1652_),
    .Y(_1745_));
 sg13g2_nand3b_1 _5257_ (.B(_2607_),
    .C(_2610_),
    .Y(_1746_),
    .A_N(_2599_));
 sg13g2_nand2b_1 _5258_ (.Y(_1747_),
    .B(_1746_),
    .A_N(_2601_));
 sg13g2_o21ai_1 _5259_ (.B1(_0641_),
    .Y(_1748_),
    .A1(net542),
    .A2(_0325_));
 sg13g2_nand2_1 _5260_ (.Y(_1749_),
    .A(_0255_),
    .B(_1748_));
 sg13g2_nand2_1 _5261_ (.Y(_1750_),
    .A(_0262_),
    .B(_1749_));
 sg13g2_a221oi_1 _5262_ (.B2(_1750_),
    .C1(_0680_),
    .B1(_0268_),
    .A1(_2562_),
    .Y(_1751_),
    .A2(_2570_));
 sg13g2_a21o_1 _5263_ (.A2(_0987_),
    .A1(_0854_),
    .B1(_1466_),
    .X(_1752_));
 sg13g2_nand2_1 _5264_ (.Y(_1753_),
    .A(_0416_),
    .B(_0418_));
 sg13g2_nor2_1 _5265_ (.A(_0411_),
    .B(_1753_),
    .Y(_1754_));
 sg13g2_mux2_1 _5266_ (.A0(_1753_),
    .A1(_1754_),
    .S(_0420_),
    .X(_1756_));
 sg13g2_a21oi_1 _5267_ (.A1(_0409_),
    .A2(_1756_),
    .Y(_1757_),
    .B1(_0328_));
 sg13g2_a21oi_1 _5268_ (.A1(net524),
    .A2(_0641_),
    .Y(_1758_),
    .B1(_0575_));
 sg13g2_or2_1 _5269_ (.X(_1759_),
    .B(_1758_),
    .A(_0620_));
 sg13g2_nand2b_1 _5270_ (.Y(_1760_),
    .B(_0825_),
    .A_N(_1036_));
 sg13g2_a22oi_1 _5271_ (.Y(_1761_),
    .B1(_0844_),
    .B2(_0713_),
    .A2(_0814_),
    .A1(net525));
 sg13g2_a22oi_1 _5272_ (.Y(_1762_),
    .B1(_0917_),
    .B2(_1760_),
    .A2(_0822_),
    .A1(net451));
 sg13g2_a21oi_1 _5273_ (.A1(net543),
    .A2(_0913_),
    .Y(_1763_),
    .B1(_0936_));
 sg13g2_o21ai_1 _5274_ (.B1(_0915_),
    .Y(_1764_),
    .A1(_1044_),
    .A2(_1763_));
 sg13g2_and4_1 _5275_ (.A(_1759_),
    .B(_1761_),
    .C(_1762_),
    .D(_1764_),
    .X(_1765_));
 sg13g2_nand3_1 _5276_ (.B(net453),
    .C(_0687_),
    .A(net490),
    .Y(_1767_));
 sg13g2_nand3_1 _5277_ (.B(_1536_),
    .C(_1767_),
    .A(_0461_),
    .Y(_1768_));
 sg13g2_nand2_1 _5278_ (.Y(_1769_),
    .A(_0614_),
    .B(_0873_));
 sg13g2_o21ai_1 _5279_ (.B1(_0908_),
    .Y(_1770_),
    .A1(_1595_),
    .A2(_1769_));
 sg13g2_a21o_1 _5280_ (.A2(_1763_),
    .A1(_1598_),
    .B1(net530),
    .X(_1771_));
 sg13g2_nand2_1 _5281_ (.Y(_1772_),
    .A(_0748_),
    .B(_0800_));
 sg13g2_a22oi_1 _5282_ (.Y(_1773_),
    .B1(_0988_),
    .B2(net531),
    .A2(net523),
    .A1(_0285_));
 sg13g2_nand3_1 _5283_ (.B(_1772_),
    .C(_1773_),
    .A(_1684_),
    .Y(_1774_));
 sg13g2_o21ai_1 _5284_ (.B1(_0805_),
    .Y(_1775_),
    .A1(net451),
    .A2(_0740_));
 sg13g2_o21ai_1 _5285_ (.B1(net489),
    .Y(_1776_),
    .A1(net519),
    .A2(net451));
 sg13g2_a221oi_1 _5286_ (.B2(_0760_),
    .C1(_1755_),
    .B1(_0759_),
    .A1(net551),
    .Y(_1778_),
    .A2(_2581_));
 sg13g2_a21oi_1 _5287_ (.A1(_1766_),
    .A2(_0761_),
    .Y(_1779_),
    .B1(net491));
 sg13g2_nor3_1 _5288_ (.A(_1081_),
    .B(_1778_),
    .C(_1779_),
    .Y(_1780_));
 sg13g2_nor4_1 _5289_ (.A(_1755_),
    .B(_2595_),
    .C(_0600_),
    .D(_1780_),
    .Y(_1781_));
 sg13g2_o21ai_1 _5290_ (.B1(_1781_),
    .Y(_1782_),
    .A1(_2583_),
    .A2(_1082_));
 sg13g2_a21oi_1 _5291_ (.A1(_0719_),
    .A2(_1782_),
    .Y(_1783_),
    .B1(_0886_));
 sg13g2_o21ai_1 _5292_ (.B1(_1496_),
    .Y(_1784_),
    .A1(net487),
    .A2(net450));
 sg13g2_a21oi_1 _5293_ (.A1(net453),
    .A2(_1784_),
    .Y(_1785_),
    .B1(_0902_));
 sg13g2_a21oi_1 _5294_ (.A1(net487),
    .A2(net455),
    .Y(_1786_),
    .B1(_0715_));
 sg13g2_nor2_1 _5295_ (.A(_0602_),
    .B(net467),
    .Y(_1787_));
 sg13g2_o21ai_1 _5296_ (.B1(_1787_),
    .Y(_1789_),
    .A1(_0687_),
    .A2(_1786_));
 sg13g2_a22oi_1 _5297_ (.Y(_1790_),
    .B1(_1789_),
    .B2(_0706_),
    .A2(_0881_),
    .A1(_0676_));
 sg13g2_nor2_1 _5298_ (.A(_0771_),
    .B(_1790_),
    .Y(_1791_));
 sg13g2_and2_1 _5299_ (.A(net447),
    .B(_1040_),
    .X(_1792_));
 sg13g2_nand2b_1 _5300_ (.Y(_1793_),
    .B(_1561_),
    .A_N(_0768_));
 sg13g2_nand2_2 _5301_ (.Y(_1794_),
    .A(_0686_),
    .B(_0772_));
 sg13g2_nand3_1 _5302_ (.B(_0775_),
    .C(_0870_),
    .A(net454),
    .Y(_1795_));
 sg13g2_nand2b_1 _5303_ (.Y(_1796_),
    .B(_0797_),
    .A_N(_0795_));
 sg13g2_o21ai_1 _5304_ (.B1(_1796_),
    .Y(_1797_),
    .A1(net489),
    .A2(net468));
 sg13g2_o21ai_1 _5305_ (.B1(_0787_),
    .Y(_1798_),
    .A1(net548),
    .A2(net481));
 sg13g2_a21oi_1 _5306_ (.A1(_1797_),
    .A2(_1798_),
    .Y(_1800_),
    .B1(net545));
 sg13g2_nand3_1 _5307_ (.B(_0806_),
    .C(_0818_),
    .A(_0753_),
    .Y(_1801_));
 sg13g2_nand3_1 _5308_ (.B(_0829_),
    .C(_0858_),
    .A(_2614_),
    .Y(_1802_));
 sg13g2_nand2_1 _5309_ (.Y(_1803_),
    .A(net526),
    .B(_0820_));
 sg13g2_nand3_1 _5310_ (.B(_1549_),
    .C(_1803_),
    .A(_0749_),
    .Y(_1804_));
 sg13g2_nor3_1 _5311_ (.A(_0329_),
    .B(_0771_),
    .C(_1786_),
    .Y(_1805_));
 sg13g2_o21ai_1 _5312_ (.B1(net522),
    .Y(_1806_),
    .A1(net545),
    .A2(net489));
 sg13g2_o21ai_1 _5313_ (.B1(_0810_),
    .Y(_1807_),
    .A1(net445),
    .A2(_1806_));
 sg13g2_nand2_1 _5314_ (.Y(_1808_),
    .A(_0647_),
    .B(_0839_));
 sg13g2_nand3_1 _5315_ (.B(_0675_),
    .C(net445),
    .A(net483),
    .Y(_1809_));
 sg13g2_o21ai_1 _5316_ (.B1(_0831_),
    .Y(_1811_),
    .A1(net525),
    .A2(_0833_));
 sg13g2_a21oi_1 _5317_ (.A1(net483),
    .A2(net520),
    .Y(_1812_),
    .B1(_0697_));
 sg13g2_nor2_1 _5318_ (.A(net546),
    .B(_2584_),
    .Y(_1813_));
 sg13g2_o21ai_1 _5319_ (.B1(_0859_),
    .Y(_1814_),
    .A1(_0733_),
    .A2(_1813_));
 sg13g2_a21oi_1 _5320_ (.A1(_0667_),
    .A2(_1053_),
    .Y(_1815_),
    .B1(_0669_));
 sg13g2_nand3_1 _5321_ (.B(_0742_),
    .C(_1055_),
    .A(net485),
    .Y(_1816_));
 sg13g2_nor3_1 _5322_ (.A(_0578_),
    .B(_0650_),
    .C(_0782_),
    .Y(_1817_));
 sg13g2_o21ai_1 _5323_ (.B1(_1809_),
    .Y(_1818_),
    .A1(_0649_),
    .A2(_0848_));
 sg13g2_a221oi_1 _5324_ (.B2(_0667_),
    .C1(_0669_),
    .B1(_1053_),
    .A1(_0655_),
    .Y(_1819_),
    .A2(_0790_));
 sg13g2_nand4_1 _5325_ (.B(_1804_),
    .C(_1816_),
    .A(_1801_),
    .Y(_1820_),
    .D(_1819_));
 sg13g2_nor4_1 _5326_ (.A(_0905_),
    .B(_0910_),
    .C(_1818_),
    .D(_1820_),
    .Y(_1822_));
 sg13g2_nand3_1 _5327_ (.B(_0709_),
    .C(_1793_),
    .A(_0688_),
    .Y(_1823_));
 sg13g2_a221oi_1 _5328_ (.B2(_0709_),
    .C1(_1774_),
    .B1(_1792_),
    .A1(_1775_),
    .Y(_1824_),
    .A2(_1776_));
 sg13g2_a221oi_1 _5329_ (.B2(_0351_),
    .C1(_1812_),
    .B1(_1662_),
    .A1(_0677_),
    .Y(_1825_),
    .A2(net464));
 sg13g2_o21ai_1 _5330_ (.B1(_1808_),
    .Y(_1826_),
    .A1(net542),
    .A2(_0920_));
 sg13g2_a221oi_1 _5331_ (.B2(net532),
    .C1(_1826_),
    .B1(_0828_),
    .A1(_0580_),
    .Y(_1827_),
    .A2(_0745_));
 sg13g2_nand4_1 _5332_ (.B(_1824_),
    .C(_1825_),
    .A(_1802_),
    .Y(_1828_),
    .D(_1827_));
 sg13g2_a221oi_1 _5333_ (.B2(_1045_),
    .C1(_1828_),
    .B1(_1771_),
    .A1(_0926_),
    .Y(_1829_),
    .A2(_1059_));
 sg13g2_nand4_1 _5334_ (.B(_1822_),
    .C(_1823_),
    .A(_1770_),
    .Y(_1830_),
    .D(_1829_));
 sg13g2_o21ai_1 _5335_ (.B1(_1795_),
    .Y(_1831_),
    .A1(_0767_),
    .A2(_1794_));
 sg13g2_a22oi_1 _5336_ (.Y(_1833_),
    .B1(_0928_),
    .B2(_0617_),
    .A2(_0721_),
    .A1(_0720_));
 sg13g2_a221oi_1 _5337_ (.B2(_1573_),
    .C1(_1817_),
    .B1(_1572_),
    .A1(_0762_),
    .Y(_1834_),
    .A2(_0764_));
 sg13g2_o21ai_1 _5338_ (.B1(_0665_),
    .Y(_1835_),
    .A1(_0748_),
    .A2(_0799_));
 sg13g2_a22oi_1 _5339_ (.Y(_1836_),
    .B1(_0741_),
    .B2(_0820_),
    .A2(_0645_),
    .A1(_0644_));
 sg13g2_a22oi_1 _5340_ (.Y(_1837_),
    .B1(_0811_),
    .B2(net531),
    .A2(_0792_),
    .A1(_0748_));
 sg13g2_nand2_1 _5341_ (.Y(_1838_),
    .A(_1836_),
    .B(_1837_));
 sg13g2_o21ai_1 _5342_ (.B1(_1814_),
    .Y(_1839_),
    .A1(_2578_),
    .A2(_2590_));
 sg13g2_nor4_2 _5343_ (.A(_1708_),
    .B(_1835_),
    .C(_1838_),
    .Y(_1840_),
    .D(_1839_));
 sg13g2_nand4_1 _5344_ (.B(_1833_),
    .C(_1834_),
    .A(_0735_),
    .Y(_1841_),
    .D(_1840_));
 sg13g2_or4_1 _5345_ (.A(_1800_),
    .B(_1805_),
    .C(_1831_),
    .D(_1841_),
    .X(_1842_));
 sg13g2_a22oi_1 _5346_ (.Y(_1844_),
    .B1(_1588_),
    .B2(_0842_),
    .A2(_1077_),
    .A1(net546));
 sg13g2_nand4_1 _5347_ (.B(_1807_),
    .C(_1811_),
    .A(_1698_),
    .Y(_1845_),
    .D(_1844_));
 sg13g2_o21ai_1 _5348_ (.B1(_1768_),
    .Y(_1846_),
    .A1(_0694_),
    .A2(_1561_));
 sg13g2_or4_1 _5349_ (.A(_1783_),
    .B(_1842_),
    .C(_1845_),
    .D(_1846_),
    .X(_1847_));
 sg13g2_nor4_2 _5350_ (.A(_1785_),
    .B(_1791_),
    .C(_1830_),
    .Y(_1848_),
    .D(_1847_));
 sg13g2_nand4_1 _5351_ (.B(_0619_),
    .C(_1765_),
    .A(_0618_),
    .Y(_1849_),
    .D(_1848_));
 sg13g2_nor3_1 _5352_ (.A(_0496_),
    .B(_1757_),
    .C(_1849_),
    .Y(_1850_));
 sg13g2_and4_1 _5353_ (.A(_1747_),
    .B(_1751_),
    .C(_1752_),
    .D(_1850_),
    .X(_1851_));
 sg13g2_a21oi_1 _5354_ (.A1(_1745_),
    .A2(_1851_),
    .Y(uo_out[6]),
    .B1(_0637_));
 sg13g2_o21ai_1 _5355_ (.B1(_2629_),
    .Y(_1852_),
    .A1(_0604_),
    .A2(_1651_));
 sg13g2_nor2_1 _5356_ (.A(_1546_),
    .B(_1671_),
    .Y(_1854_));
 sg13g2_nand3_1 _5357_ (.B(_0409_),
    .C(_1756_),
    .A(_0330_),
    .Y(_1855_));
 sg13g2_nand2b_1 _5358_ (.Y(_1856_),
    .B(_0645_),
    .A_N(_0644_));
 sg13g2_o21ai_1 _5359_ (.B1(_1856_),
    .Y(_1857_),
    .A1(_0699_),
    .A2(_0819_));
 sg13g2_a221oi_1 _5360_ (.B2(_1070_),
    .C1(_1857_),
    .B1(net464),
    .A1(_0748_),
    .Y(_1858_),
    .A2(_0810_));
 sg13g2_nand2_1 _5361_ (.Y(_1859_),
    .A(_0675_),
    .B(_0733_));
 sg13g2_a21oi_1 _5362_ (.A1(net483),
    .A2(net451),
    .Y(_1860_),
    .B1(_0805_));
 sg13g2_a21oi_1 _5363_ (.A1(_0646_),
    .A2(_0839_),
    .Y(_1861_),
    .B1(_1860_));
 sg13g2_nand4_1 _5364_ (.B(_1858_),
    .C(_1859_),
    .A(_1794_),
    .Y(_1862_),
    .D(_1861_));
 sg13g2_a21oi_1 _5365_ (.A1(net492),
    .A2(net464),
    .Y(_1863_),
    .B1(_0682_));
 sg13g2_a221oi_1 _5366_ (.B2(_0921_),
    .C1(_1863_),
    .B1(_0855_),
    .A1(_0649_),
    .Y(_1865_),
    .A2(_0829_));
 sg13g2_nand3_1 _5367_ (.B(net468),
    .C(_0828_),
    .A(net522),
    .Y(_1866_));
 sg13g2_nand3_1 _5368_ (.B(_0498_),
    .C(_0858_),
    .A(_0266_),
    .Y(_1867_));
 sg13g2_a22oi_1 _5369_ (.Y(_1868_),
    .B1(_1071_),
    .B2(_0650_),
    .A2(_0664_),
    .A1(_0661_));
 sg13g2_nand4_1 _5370_ (.B(_1866_),
    .C(_1867_),
    .A(_1865_),
    .Y(_1869_),
    .D(_1868_));
 sg13g2_nor4_1 _5371_ (.A(_0676_),
    .B(_0764_),
    .C(_0908_),
    .D(_0942_),
    .Y(_1870_));
 sg13g2_nor2_1 _5372_ (.A(_0739_),
    .B(_0831_),
    .Y(_1871_));
 sg13g2_a21oi_1 _5373_ (.A1(net456),
    .A2(_0729_),
    .Y(_1872_),
    .B1(_1075_));
 sg13g2_nand4_1 _5374_ (.B(_1870_),
    .C(_1871_),
    .A(_0406_),
    .Y(_1873_),
    .D(_1872_));
 sg13g2_a21oi_1 _5375_ (.A1(_0749_),
    .A2(_0752_),
    .Y(_1874_),
    .B1(_1579_));
 sg13g2_a22oi_1 _5376_ (.Y(_1876_),
    .B1(net464),
    .B2(_0677_),
    .A2(_0781_),
    .A1(_0579_));
 sg13g2_nor2_1 _5377_ (.A(_2579_),
    .B(_1062_),
    .Y(_1877_));
 sg13g2_nand4_1 _5378_ (.B(_1874_),
    .C(_1876_),
    .A(_1104_),
    .Y(_1878_),
    .D(_1877_));
 sg13g2_or4_1 _5379_ (.A(_1862_),
    .B(_1869_),
    .C(_1873_),
    .D(_1878_),
    .X(_1879_));
 sg13g2_a21oi_1 _5380_ (.A1(net457),
    .A2(_0691_),
    .Y(_1880_),
    .B1(net470));
 sg13g2_nand3_1 _5381_ (.B(net453),
    .C(_1880_),
    .A(_0603_),
    .Y(_1881_));
 sg13g2_nand3_1 _5382_ (.B(_0614_),
    .C(_0910_),
    .A(net455),
    .Y(_1882_));
 sg13g2_o21ai_1 _5383_ (.B1(_0870_),
    .Y(_1883_),
    .A1(net488),
    .A2(_0603_));
 sg13g2_nand3_1 _5384_ (.B(_1882_),
    .C(_1883_),
    .A(_1881_),
    .Y(_1884_));
 sg13g2_a21oi_1 _5385_ (.A1(_0708_),
    .A2(_0900_),
    .Y(_1885_),
    .B1(_1774_));
 sg13g2_a22oi_1 _5386_ (.Y(_1887_),
    .B1(_1077_),
    .B2(_1317_),
    .A2(_0787_),
    .A1(_0784_));
 sg13g2_nand3_1 _5387_ (.B(_0688_),
    .C(_0770_),
    .A(_0603_),
    .Y(_1888_));
 sg13g2_nand3_1 _5388_ (.B(_1887_),
    .C(_1888_),
    .A(_1885_),
    .Y(_1889_));
 sg13g2_nor2_1 _5389_ (.A(_0720_),
    .B(_0904_),
    .Y(_1890_));
 sg13g2_a221oi_1 _5390_ (.B2(_1673_),
    .C1(_1890_),
    .B1(_1787_),
    .A1(_0461_),
    .Y(_1891_),
    .A2(_1697_));
 sg13g2_o21ai_1 _5391_ (.B1(net521),
    .Y(_1892_),
    .A1(net481),
    .A2(_0658_));
 sg13g2_a22oi_1 _5392_ (.Y(_1893_),
    .B1(_1892_),
    .B2(_0742_),
    .A2(_1040_),
    .A1(_0875_));
 sg13g2_a221oi_1 _5393_ (.B2(_0527_),
    .C1(_0860_),
    .B1(_2603_),
    .A1(net539),
    .Y(_1894_),
    .A2(_2584_));
 sg13g2_a21oi_1 _5394_ (.A1(_0741_),
    .A2(_0807_),
    .Y(_1895_),
    .B1(_1894_));
 sg13g2_nand2_1 _5395_ (.Y(_1896_),
    .A(_1893_),
    .B(_1895_));
 sg13g2_o21ai_1 _5396_ (.B1(_1815_),
    .Y(_1898_),
    .A1(_0789_),
    .A2(_1055_));
 sg13g2_nor4_1 _5397_ (.A(_1057_),
    .B(_1705_),
    .C(_1896_),
    .D(_1898_),
    .Y(_1899_));
 sg13g2_or2_1 _5398_ (.X(_1900_),
    .B(_1595_),
    .A(_1594_));
 sg13g2_nand4_1 _5399_ (.B(_1891_),
    .C(_1899_),
    .A(_1700_),
    .Y(_1901_),
    .D(_1900_));
 sg13g2_nor4_1 _5400_ (.A(_1879_),
    .B(_1884_),
    .C(_1889_),
    .D(_1901_),
    .Y(_1902_));
 sg13g2_a21oi_1 _5401_ (.A1(_0913_),
    .A2(_1675_),
    .Y(_1903_),
    .B1(_0936_));
 sg13g2_o21ai_1 _5402_ (.B1(_1045_),
    .Y(_1904_),
    .A1(net530),
    .A2(_1903_));
 sg13g2_or3_1 _5403_ (.A(_2626_),
    .B(net469),
    .C(_1049_),
    .X(_1905_));
 sg13g2_nand4_1 _5404_ (.B(_1902_),
    .C(_1904_),
    .A(_1126_),
    .Y(_1906_),
    .D(_1905_));
 sg13g2_nor2_1 _5405_ (.A(_1127_),
    .B(_1906_),
    .Y(_1907_));
 sg13g2_and3_1 _5406_ (.X(_1909_),
    .A(_1765_),
    .B(_1855_),
    .C(_1907_));
 sg13g2_o21ai_1 _5407_ (.B1(_1909_),
    .Y(_1910_),
    .A1(_1466_),
    .A2(_1854_));
 sg13g2_and2_1 _5408_ (.A(_1751_),
    .B(_1852_),
    .X(_1911_));
 sg13g2_nor2_1 _5409_ (.A(_1000_),
    .B(_1910_),
    .Y(_1912_));
 sg13g2_a21oi_1 _5410_ (.A1(_1911_),
    .A2(_1912_),
    .Y(uo_out[2]),
    .B1(_0637_));
 sg13g2_nand3_1 _5411_ (.B(_2670_),
    .C(_0359_),
    .A(_0648_),
    .Y(_1913_));
 sg13g2_nor3_2 _5412_ (.A(net552),
    .B(net551),
    .C(_1913_),
    .Y(_1914_));
 sg13g2_nor2_2 _5413_ (.A(_0043_),
    .B(_1914_),
    .Y(_1915_));
 sg13g2_nand2b_2 _5414_ (.Y(_1916_),
    .B(net656),
    .A_N(_1914_));
 sg13g2_nor2_1 _5415_ (.A(net647),
    .B(_1916_),
    .Y(_0000_));
 sg13g2_nor2_1 _5416_ (.A(_1021_),
    .B(_1916_),
    .Y(_0001_));
 sg13g2_and2_1 _5417_ (.A(_2680_),
    .B(_1915_),
    .X(_0002_));
 sg13g2_nor2_1 _5418_ (.A(_2673_),
    .B(_1916_),
    .Y(_0003_));
 sg13g2_nor2_1 _5419_ (.A(_0043_),
    .B(_1140_),
    .Y(_0004_));
 sg13g2_nor2_2 _5420_ (.A(_2557_),
    .B(_2671_),
    .Y(_1918_));
 sg13g2_a21oi_1 _5421_ (.A1(net632),
    .A2(_2670_),
    .Y(_1919_),
    .B1(net631));
 sg13g2_nor3_1 _5422_ (.A(_1916_),
    .B(_1918_),
    .C(net69),
    .Y(_0005_));
 sg13g2_o21ai_1 _5423_ (.B1(_1915_),
    .Y(_1920_),
    .A1(net625),
    .A2(_1918_));
 sg13g2_a21oi_1 _5424_ (.A1(net625),
    .A2(_1918_),
    .Y(_0006_),
    .B1(_1920_));
 sg13g2_a21oi_1 _5425_ (.A1(net625),
    .A2(_1918_),
    .Y(_1921_),
    .B1(net620));
 sg13g2_nor3_1 _5426_ (.A(_2553_),
    .B(_2557_),
    .C(_2671_),
    .Y(_1923_));
 sg13g2_nor3_1 _5427_ (.A(_1916_),
    .B(_1921_),
    .C(_1923_),
    .Y(_0007_));
 sg13g2_nor2_1 _5428_ (.A(net615),
    .B(_1923_),
    .Y(_1924_));
 sg13g2_and2_1 _5429_ (.A(net615),
    .B(_1923_),
    .X(_1925_));
 sg13g2_nor3_1 _5430_ (.A(_1916_),
    .B(_1924_),
    .C(_1925_),
    .Y(_0008_));
 sg13g2_xnor2_1 _5431_ (.Y(_1926_),
    .A(net610),
    .B(_1925_));
 sg13g2_nor2_1 _5432_ (.A(_1916_),
    .B(_1926_),
    .Y(_0009_));
 sg13g2_a21o_1 _5433_ (.A2(_2657_),
    .A1(net3),
    .B1(net5),
    .X(_0010_));
 sg13g2_or2_1 _5434_ (.X(_0011_),
    .B(net4),
    .A(net5));
 sg13g2_or3_1 _5435_ (.A(net3),
    .B(net2),
    .C(_0011_),
    .X(_0012_));
 sg13g2_nand3_1 _5436_ (.B(net655),
    .C(_2620_),
    .A(net608),
    .Y(_1928_));
 sg13g2_a221oi_1 _5437_ (.B2(_2556_),
    .C1(_1928_),
    .B1(_2552_),
    .A1(net556),
    .Y(_0013_),
    .A2(_0912_));
 sg13g2_nand2b_1 _5438_ (.Y(_1929_),
    .B(net656),
    .A_N(net55));
 sg13g2_nor4_2 _5439_ (.A(_0593_),
    .B(_0823_),
    .C(_0911_),
    .Y(_0014_),
    .D(_1929_));
 sg13g2_nand2_1 _5440_ (.Y(_1930_),
    .A(\hvsync_gen.vpos[9] ),
    .B(_1218_));
 sg13g2_or4_1 _5441_ (.A(net544),
    .B(_2447_),
    .C(_0606_),
    .D(_1930_),
    .X(_1931_));
 sg13g2_a21o_1 _5442_ (.A2(_1931_),
    .A1(_1914_),
    .B1(net601),
    .X(_1932_));
 sg13g2_nand2_1 _5443_ (.Y(_1933_),
    .A(net602),
    .B(_1914_));
 sg13g2_and3_1 _5444_ (.X(_0015_),
    .A(net656),
    .B(_1932_),
    .C(_1933_));
 sg13g2_a221oi_1 _5445_ (.B2(_2624_),
    .C1(_0043_),
    .B1(_1933_),
    .A1(_0425_),
    .Y(_0016_),
    .A2(_1914_));
 sg13g2_nand2_1 _5446_ (.Y(_1935_),
    .A(net595),
    .B(_1915_));
 sg13g2_xnor2_1 _5447_ (.Y(_1936_),
    .A(_2613_),
    .B(_0426_));
 sg13g2_nand3_1 _5448_ (.B(_1914_),
    .C(_1931_),
    .A(net656),
    .Y(_1937_));
 sg13g2_o21ai_1 _5449_ (.B1(_1935_),
    .Y(_0017_),
    .A1(_1936_),
    .A2(_1937_));
 sg13g2_a21oi_1 _5450_ (.A1(net597),
    .A2(_0425_),
    .Y(_1938_),
    .B1(net592));
 sg13g2_nor2_1 _5451_ (.A(_2447_),
    .B(_0426_),
    .Y(_1939_));
 sg13g2_or3_1 _5452_ (.A(_1937_),
    .B(_1938_),
    .C(_1939_),
    .X(_1940_));
 sg13g2_o21ai_1 _5453_ (.B1(_1940_),
    .Y(_0018_),
    .A1(net561),
    .A2(_1916_));
 sg13g2_and2_1 _5454_ (.A(_1914_),
    .B(_1939_),
    .X(_1941_));
 sg13g2_nand2_1 _5455_ (.Y(_1942_),
    .A(_1914_),
    .B(_1939_));
 sg13g2_nand2_1 _5456_ (.Y(_1944_),
    .A(net587),
    .B(_1941_));
 sg13g2_nand2_1 _5457_ (.Y(_1945_),
    .A(net656),
    .B(_1944_));
 sg13g2_a21oi_1 _5458_ (.A1(_2591_),
    .A2(_1942_),
    .Y(_0019_),
    .B1(_1945_));
 sg13g2_a221oi_1 _5459_ (.B2(_2580_),
    .C1(_0043_),
    .B1(_1944_),
    .A1(_1131_),
    .Y(_0020_),
    .A2(_1941_));
 sg13g2_a21oi_1 _5460_ (.A1(_1131_),
    .A2(_1941_),
    .Y(_1946_),
    .B1(net579));
 sg13g2_nor2_1 _5461_ (.A(_1493_),
    .B(_1942_),
    .Y(_1947_));
 sg13g2_nor3_1 _5462_ (.A(_0043_),
    .B(_1946_),
    .C(_1947_),
    .Y(_0021_));
 sg13g2_o21ai_1 _5463_ (.B1(net656),
    .Y(_1948_),
    .A1(net572),
    .A2(_1947_));
 sg13g2_a21oi_1 _5464_ (.A1(_1163_),
    .A2(_1941_),
    .Y(_0022_),
    .B1(_1948_));
 sg13g2_a21oi_1 _5465_ (.A1(_1163_),
    .A2(_1941_),
    .Y(_1949_),
    .B1(net566));
 sg13g2_nor2_1 _5466_ (.A(_0593_),
    .B(_1944_),
    .Y(_1951_));
 sg13g2_nor3_1 _5467_ (.A(_0043_),
    .B(_1949_),
    .C(_1951_),
    .Y(_0023_));
 sg13g2_nand2_1 _5468_ (.Y(_1952_),
    .A(net55),
    .B(_1915_));
 sg13g2_nand3_1 _5469_ (.B(_1163_),
    .C(_1939_),
    .A(net566),
    .Y(_1953_));
 sg13g2_xor2_1 _5470_ (.B(_1953_),
    .A(net55),
    .X(_1954_));
 sg13g2_o21ai_1 _5471_ (.B1(_1952_),
    .Y(_0024_),
    .A1(_1937_),
    .A2(_1954_));
 sg13g2_or2_1 _5472_ (.X(_1955_),
    .B(_0012_),
    .A(_0032_));
 sg13g2_a21oi_1 _5473_ (.A1(\reset_latch[1] ),
    .A2(\reset_latch[0] ),
    .Y(_1956_),
    .B1(net517));
 sg13g2_a21o_2 _5474_ (.A2(\reset_latch[0] ),
    .A1(\reset_latch[1] ),
    .B1(net517),
    .X(_1957_));
 sg13g2_nand2_1 _5475_ (.Y(_1958_),
    .A(\reset_latch[2] ),
    .B(\reset_latch[0] ));
 sg13g2_nor2_2 _5476_ (.A(\reset_latch[1] ),
    .B(_1958_),
    .Y(_1960_));
 sg13g2_or2_1 _5477_ (.X(_1961_),
    .B(_1958_),
    .A(\reset_latch[1] ));
 sg13g2_nand3b_1 _5478_ (.B(\reset_latch[1] ),
    .C(\reset_latch[2] ),
    .Y(_1962_),
    .A_N(\reset_latch[0] ));
 sg13g2_nor2_1 _5479_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .Y(_1963_));
 sg13g2_o21ai_1 _5480_ (.B1(\counter[2] ),
    .Y(_1964_),
    .A1(\counter[1] ),
    .A2(\counter[0] ));
 sg13g2_nand2_1 _5481_ (.Y(_1965_),
    .A(_0054_),
    .B(_1964_));
 sg13g2_a21oi_1 _5482_ (.A1(\counter[4] ),
    .A2(_1965_),
    .Y(_1966_),
    .B1(\counter[5] ));
 sg13g2_nand2b_1 _5483_ (.Y(_1967_),
    .B(net56),
    .A_N(_1966_));
 sg13g2_nor2b_2 _5484_ (.A(net540),
    .B_N(_1967_),
    .Y(_1968_));
 sg13g2_nor2_1 _5485_ (.A(_1960_),
    .B(_1968_),
    .Y(_1969_));
 sg13g2_nand3_1 _5486_ (.B(_1961_),
    .C(net540),
    .A(net6),
    .Y(_1971_));
 sg13g2_o21ai_1 _5487_ (.B1(_1971_),
    .Y(_1972_),
    .A1(net62),
    .A2(_1969_));
 sg13g2_a22oi_1 _5488_ (.Y(_1973_),
    .B1(_1956_),
    .B2(_1972_),
    .A2(net517),
    .A1(net62));
 sg13g2_inv_1 _5489_ (.Y(_0025_),
    .A(net63));
 sg13g2_and2_1 _5490_ (.A(\counter[1] ),
    .B(\counter[0] ),
    .X(_1974_));
 sg13g2_nor2_1 _5491_ (.A(_1963_),
    .B(_1974_),
    .Y(_1975_));
 sg13g2_nand2b_2 _5492_ (.Y(_1976_),
    .B(_1963_),
    .A_N(\counter[2] ));
 sg13g2_nor2_1 _5493_ (.A(\counter[3] ),
    .B(_1976_),
    .Y(_1977_));
 sg13g2_nor3_1 _5494_ (.A(\counter[4] ),
    .B(\counter[3] ),
    .C(_1976_),
    .Y(_1978_));
 sg13g2_or2_1 _5495_ (.X(_1979_),
    .B(net56),
    .A(\counter[5] ));
 sg13g2_nand2b_1 _5496_ (.Y(_1981_),
    .B(_1978_),
    .A_N(\counter[5] ));
 sg13g2_o21ai_1 _5497_ (.B1(_1960_),
    .Y(_1982_),
    .A1(\counter[6] ),
    .A2(_1981_));
 sg13g2_nor2_1 _5498_ (.A(_1975_),
    .B(_1982_),
    .Y(_1983_));
 sg13g2_a21oi_1 _5499_ (.A1(net7),
    .A2(_1961_),
    .Y(_1984_),
    .B1(_1983_));
 sg13g2_a21o_1 _5500_ (.A2(_1975_),
    .A1(_1967_),
    .B1(net540),
    .X(_1985_));
 sg13g2_a21oi_1 _5501_ (.A1(net540),
    .A2(_1984_),
    .Y(_1986_),
    .B1(_1957_));
 sg13g2_a22oi_1 _5502_ (.Y(_1987_),
    .B1(_1985_),
    .B2(_1986_),
    .A2(net517),
    .A1(net58));
 sg13g2_inv_1 _5503_ (.Y(_0026_),
    .A(net59));
 sg13g2_nand2_1 _5504_ (.Y(_1988_),
    .A(\counter[2] ),
    .B(_1974_));
 sg13g2_xor2_1 _5505_ (.B(_1974_),
    .A(\counter[2] ),
    .X(_1989_));
 sg13g2_nand3_1 _5506_ (.B(_1961_),
    .C(_1962_),
    .A(net8),
    .Y(_1991_));
 sg13g2_nand2_1 _5507_ (.Y(_1992_),
    .A(_1964_),
    .B(_1976_));
 sg13g2_a22oi_1 _5508_ (.Y(_1993_),
    .B1(_1992_),
    .B2(_1960_),
    .A2(_1989_),
    .A1(_1968_));
 sg13g2_a21oi_1 _5509_ (.A1(_1991_),
    .A2(_1993_),
    .Y(_1994_),
    .B1(_1957_));
 sg13g2_a21o_1 _5510_ (.A2(_1955_),
    .A1(net60),
    .B1(_1994_),
    .X(_0027_));
 sg13g2_nand2_1 _5511_ (.Y(_1995_),
    .A(net51),
    .B(net517));
 sg13g2_xnor2_1 _5512_ (.Y(_1996_),
    .A(_0054_),
    .B(_1976_));
 sg13g2_nand2_1 _5513_ (.Y(_1997_),
    .A(net9),
    .B(_1961_));
 sg13g2_o21ai_1 _5514_ (.B1(_1997_),
    .Y(_1998_),
    .A1(_1982_),
    .A2(_1996_));
 sg13g2_nor2_1 _5515_ (.A(_0054_),
    .B(_1988_),
    .Y(_1999_));
 sg13g2_xnor2_1 _5516_ (.Y(_2001_),
    .A(net51),
    .B(_1988_));
 sg13g2_a22oi_1 _5517_ (.Y(_2002_),
    .B1(_2001_),
    .B2(_1968_),
    .A2(_1998_),
    .A1(net540));
 sg13g2_o21ai_1 _5518_ (.B1(_1995_),
    .Y(_0028_),
    .A1(_1957_),
    .A2(_2002_));
 sg13g2_nand2_1 _5519_ (.Y(_2003_),
    .A(\counter[4] ),
    .B(_1999_));
 sg13g2_xor2_1 _5520_ (.B(_1999_),
    .A(\counter[4] ),
    .X(_2004_));
 sg13g2_xor2_1 _5521_ (.B(_1977_),
    .A(net65),
    .X(_2005_));
 sg13g2_nand3_1 _5522_ (.B(_1961_),
    .C(net540),
    .A(net10),
    .Y(_2006_));
 sg13g2_a22oi_1 _5523_ (.Y(_2007_),
    .B1(_2005_),
    .B2(_1960_),
    .A2(_2004_),
    .A1(_1968_));
 sg13g2_a21oi_1 _5524_ (.A1(_2006_),
    .A2(_2007_),
    .Y(_2008_),
    .B1(_1957_));
 sg13g2_a21o_1 _5525_ (.A2(net517),
    .A1(net65),
    .B1(_2008_),
    .X(_0029_));
 sg13g2_nand2_1 _5526_ (.Y(_2010_),
    .A(net53),
    .B(net517));
 sg13g2_xnor2_1 _5527_ (.Y(_2011_),
    .A(\counter[5] ),
    .B(_1978_));
 sg13g2_nand2_1 _5528_ (.Y(_2012_),
    .A(net11),
    .B(_1961_));
 sg13g2_o21ai_1 _5529_ (.B1(_2012_),
    .Y(_2013_),
    .A1(_1982_),
    .A2(_2011_));
 sg13g2_xnor2_1 _5530_ (.Y(_2014_),
    .A(net53),
    .B(_2003_));
 sg13g2_a22oi_1 _5531_ (.Y(_2015_),
    .B1(_2014_),
    .B2(_1968_),
    .A2(_2013_),
    .A1(net540));
 sg13g2_o21ai_1 _5532_ (.B1(_2010_),
    .Y(_0030_),
    .A1(_1957_),
    .A2(_2015_));
 sg13g2_nand2b_1 _5533_ (.Y(_2016_),
    .B(_2003_),
    .A_N(_1966_));
 sg13g2_nand3_1 _5534_ (.B(_1979_),
    .C(_2016_),
    .A(_1968_),
    .Y(_2017_));
 sg13g2_a21oi_1 _5535_ (.A1(net56),
    .A2(_1981_),
    .Y(_2018_),
    .B1(_1982_));
 sg13g2_a21oi_1 _5536_ (.A1(net12),
    .A2(net540),
    .Y(_2020_),
    .B1(_1960_));
 sg13g2_o21ai_1 _5537_ (.B1(_2017_),
    .Y(_2021_),
    .A1(_2018_),
    .A2(_2020_));
 sg13g2_a22oi_1 _5538_ (.Y(_2022_),
    .B1(_1956_),
    .B2(_2021_),
    .A2(net517),
    .A1(net56));
 sg13g2_inv_1 _5539_ (.Y(_0031_),
    .A(net57));
 sg13g2_dfrbpq_2 _5540_ (.RESET_B(net40),
    .D(_0000_),
    .Q(\flag.flag_abrosexual_inst.pix_x[0] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _5541_ (.RESET_B(net32),
    .D(_0001_),
    .Q(\flag.flag_abrosexual_inst.pix_x[1] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _5542_ (.RESET_B(net31),
    .D(_0002_),
    .Q(\flag.flag_abrosexual_inst.pix_x[2] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _5543_ (.RESET_B(net30),
    .D(_0003_),
    .Q(\flag.flag_abrosexual_inst.pix_x[3] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _5544_ (.RESET_B(net29),
    .D(_0004_),
    .Q(\flag.flag_abrosexual_inst.pix_x[4] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _5545_ (.RESET_B(net50),
    .D(_0005_),
    .Q(\flag.flag_abrosexual_inst.pix_x[5] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _5546_ (.RESET_B(net49),
    .D(_0006_),
    .Q(\flag.flag_abrosexual_inst.pix_x[6] ),
    .CLK(clknet_3_1__leaf_clk));
 sg13g2_dfrbpq_1 _5547_ (.RESET_B(net48),
    .D(_0007_),
    .Q(\flag.flag_abrosexual_inst.pix_x[7] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _5548_ (.RESET_B(net47),
    .D(_0008_),
    .Q(\flag.flag_abrosexual_inst.pix_x[8] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_1 _5549_ (.RESET_B(net46),
    .D(_0009_),
    .Q(\flag.flag_abrosexual_inst.pix_x[9] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_2 _5550_ (.RESET_B(net654),
    .D(_0010_),
    .Q(\reset_latch[0] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _5551_ (.RESET_B(net654),
    .D(_0011_),
    .Q(\reset_latch[1] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _5552_ (.RESET_B(net654),
    .D(_0012_),
    .Q(\reset_latch[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_1 _5553_ (.RESET_B(net45),
    .D(_0013_),
    .Q(hsync),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _5554_ (.RESET_B(net44),
    .D(net71),
    .Q(\hvsync_gen.vsync ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_1 _5555_ (.RESET_B(net43),
    .D(_0015_),
    .Q(\flag.flag_abrosexual_inst.pix_y[0] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _5556_ (.RESET_B(net41),
    .D(net79),
    .Q(\flag.flag_abrosexual_inst.pix_y[1] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_1 _5557_ (.RESET_B(net39),
    .D(_0017_),
    .Q(\flag.flag_abrosexual_inst.pix_y[2] ),
    .CLK(clknet_3_3__leaf_clk));
 sg13g2_dfrbpq_1 _5558_ (.RESET_B(net38),
    .D(_0018_),
    .Q(\flag.flag_abrosexual_inst.pix_y[3] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _5559_ (.RESET_B(net37),
    .D(_0019_),
    .Q(\flag.flag_abrosexual_inst.pix_y[4] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _5560_ (.RESET_B(net36),
    .D(_0020_),
    .Q(\flag.flag_abrosexual_inst.pix_y[5] ),
    .CLK(clknet_3_0__leaf_clk));
 sg13g2_dfrbpq_2 _5561_ (.RESET_B(net35),
    .D(_0021_),
    .Q(\flag.flag_abrosexual_inst.pix_y[6] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _5562_ (.RESET_B(net34),
    .D(_0022_),
    .Q(\flag.flag_abrosexual_inst.pix_y[7] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _5563_ (.RESET_B(net33),
    .D(_0023_),
    .Q(\flag.flag_abrosexual_inst.pix_y[8] ),
    .CLK(clknet_3_4__leaf_clk));
 sg13g2_dfrbpq_2 _5564_ (.RESET_B(net42),
    .D(_0024_),
    .Q(\hvsync_gen.vpos[9] ),
    .CLK(clknet_3_2__leaf_clk));
 sg13g2_dfrbpq_2 _5565_ (.RESET_B(net654),
    .D(_0025_),
    .Q(\counter[0] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _5566_ (.RESET_B(net654),
    .D(_0026_),
    .Q(\counter[1] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _5567_ (.RESET_B(net655),
    .D(net61),
    .Q(\counter[2] ),
    .CLK(clknet_3_7__leaf_clk));
 sg13g2_dfrbpq_2 _5568_ (.RESET_B(net655),
    .D(net52),
    .Q(\counter[3] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _5569_ (.RESET_B(net654),
    .D(net66),
    .Q(\counter[4] ),
    .CLK(clknet_3_6__leaf_clk));
 sg13g2_dfrbpq_2 _5570_ (.RESET_B(net654),
    .D(net54),
    .Q(\counter[5] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_dfrbpq_2 _5571_ (.RESET_B(net654),
    .D(_0031_),
    .Q(\counter[6] ),
    .CLK(clknet_3_5__leaf_clk));
 sg13g2_tiehi _5543__30 (.L_HI(net30));
 sg13g2_tiehi _5542__31 (.L_HI(net31));
 sg13g2_tiehi _5541__32 (.L_HI(net32));
 sg13g2_tiehi _5563__33 (.L_HI(net33));
 sg13g2_tiehi _5562__34 (.L_HI(net34));
 sg13g2_tiehi _5561__35 (.L_HI(net35));
 sg13g2_tiehi _5560__36 (.L_HI(net36));
 sg13g2_tiehi _5559__37 (.L_HI(net37));
 sg13g2_tiehi _5558__38 (.L_HI(net38));
 sg13g2_tiehi _5557__39 (.L_HI(net39));
 sg13g2_tiehi _5540__40 (.L_HI(net40));
 sg13g2_tiehi _5556__41 (.L_HI(net41));
 sg13g2_tiehi _5564__42 (.L_HI(net42));
 sg13g2_tiehi _5555__43 (.L_HI(net43));
 sg13g2_tiehi _5554__44 (.L_HI(net44));
 sg13g2_tiehi _5553__45 (.L_HI(net45));
 sg13g2_tiehi _5549__46 (.L_HI(net46));
 sg13g2_tiehi _5548__47 (.L_HI(net47));
 sg13g2_tiehi _5547__48 (.L_HI(net48));
 sg13g2_tiehi _5546__49 (.L_HI(net49));
 sg13g2_tiehi _5545__50 (.L_HI(net50));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_14 (.L_LO(net14));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_15 (.L_LO(net15));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_16 (.L_LO(net16));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_17 (.L_LO(net17));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_18 (.L_LO(net18));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_19 (.L_LO(net19));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_20 (.L_LO(net20));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_21 (.L_LO(net21));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_22 (.L_LO(net22));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_23 (.L_LO(net23));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_24 (.L_LO(net24));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_25 (.L_LO(net25));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_26 (.L_LO(net26));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_27 (.L_LO(net27));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_28 (.L_LO(net28));
 sg13g2_tiehi _5544__29 (.L_HI(net29));
 sg13g2_buf_1 _5610_ (.A(\hvsync_gen.vsync ),
    .X(uo_out[3]));
 sg13g2_buf_1 _5611_ (.A(hsync),
    .X(uo_out[7]));
 sg13g2_buf_8 fanout444 (.A(_0718_),
    .X(net444));
 sg13g2_buf_8 fanout445 (.A(_0746_),
    .X(net445));
 sg13g2_buf_8 fanout446 (.A(_0713_),
    .X(net446));
 sg13g2_buf_8 fanout447 (.A(_0603_),
    .X(net447));
 sg13g2_buf_8 fanout448 (.A(_1188_),
    .X(net448));
 sg13g2_buf_8 fanout449 (.A(_1179_),
    .X(net449));
 sg13g2_buf_8 fanout450 (.A(_0686_),
    .X(net450));
 sg13g2_buf_8 fanout451 (.A(_0660_),
    .X(net451));
 sg13g2_buf_8 fanout452 (.A(_0610_),
    .X(net452));
 sg13g2_buf_8 fanout453 (.A(_0609_),
    .X(net453));
 sg13g2_buf_8 fanout454 (.A(_0609_),
    .X(net454));
 sg13g2_buf_8 fanout455 (.A(_0601_),
    .X(net455));
 sg13g2_buf_2 fanout456 (.A(_0601_),
    .X(net456));
 sg13g2_buf_8 fanout457 (.A(_0589_),
    .X(net457));
 sg13g2_buf_8 fanout458 (.A(_2695_),
    .X(net458));
 sg13g2_buf_8 fanout459 (.A(_2676_),
    .X(net459));
 sg13g2_buf_8 fanout460 (.A(_2041_),
    .X(net460));
 sg13g2_buf_8 fanout461 (.A(_1799_),
    .X(net461));
 sg13g2_buf_8 fanout462 (.A(_1361_),
    .X(net462));
 sg13g2_buf_1 fanout463 (.A(_1361_),
    .X(net463));
 sg13g2_buf_8 fanout464 (.A(_0854_),
    .X(net464));
 sg13g2_buf_8 fanout465 (.A(net466),
    .X(net465));
 sg13g2_buf_8 fanout466 (.A(_0674_),
    .X(net466));
 sg13g2_buf_8 fanout467 (.A(_0613_),
    .X(net467));
 sg13g2_buf_8 fanout468 (.A(_0579_),
    .X(net468));
 sg13g2_buf_8 fanout469 (.A(net470),
    .X(net469));
 sg13g2_buf_8 fanout470 (.A(net471),
    .X(net470));
 sg13g2_buf_8 fanout471 (.A(_0499_),
    .X(net471));
 sg13g2_buf_8 fanout472 (.A(net474),
    .X(net472));
 sg13g2_buf_8 fanout473 (.A(net474),
    .X(net473));
 sg13g2_buf_8 fanout474 (.A(_0265_),
    .X(net474));
 sg13g2_buf_8 fanout475 (.A(_0239_),
    .X(net475));
 sg13g2_buf_8 fanout476 (.A(_0224_),
    .X(net476));
 sg13g2_buf_8 fanout477 (.A(_2628_),
    .X(net477));
 sg13g2_buf_8 fanout478 (.A(net479),
    .X(net478));
 sg13g2_buf_8 fanout479 (.A(_2628_),
    .X(net479));
 sg13g2_buf_8 fanout480 (.A(net482),
    .X(net480));
 sg13g2_buf_1 fanout481 (.A(net482),
    .X(net481));
 sg13g2_buf_8 fanout482 (.A(_2586_),
    .X(net482));
 sg13g2_buf_8 fanout483 (.A(net485),
    .X(net483));
 sg13g2_buf_1 fanout484 (.A(net485),
    .X(net484));
 sg13g2_buf_8 fanout485 (.A(net486),
    .X(net485));
 sg13g2_buf_2 fanout486 (.A(_2586_),
    .X(net486));
 sg13g2_buf_8 fanout487 (.A(net488),
    .X(net487));
 sg13g2_buf_2 fanout488 (.A(net490),
    .X(net488));
 sg13g2_buf_8 fanout489 (.A(net490),
    .X(net489));
 sg13g2_buf_8 fanout490 (.A(_2585_),
    .X(net490));
 sg13g2_buf_8 fanout491 (.A(net494),
    .X(net491));
 sg13g2_buf_8 fanout492 (.A(net494),
    .X(net492));
 sg13g2_buf_1 fanout493 (.A(net494),
    .X(net493));
 sg13g2_buf_8 fanout494 (.A(_2585_),
    .X(net494));
 sg13g2_buf_8 fanout495 (.A(_2566_),
    .X(net495));
 sg13g2_buf_8 fanout496 (.A(_2566_),
    .X(net496));
 sg13g2_buf_8 fanout497 (.A(net498),
    .X(net497));
 sg13g2_buf_8 fanout498 (.A(_2330_),
    .X(net498));
 sg13g2_buf_8 fanout499 (.A(net500),
    .X(net499));
 sg13g2_buf_8 fanout500 (.A(_2048_),
    .X(net500));
 sg13g2_buf_8 fanout501 (.A(net502),
    .X(net501));
 sg13g2_buf_8 fanout502 (.A(_2040_),
    .X(net502));
 sg13g2_buf_8 fanout503 (.A(net504),
    .X(net503));
 sg13g2_buf_8 fanout504 (.A(_2034_),
    .X(net504));
 sg13g2_buf_8 fanout505 (.A(_2026_),
    .X(net505));
 sg13g2_buf_8 fanout506 (.A(_2026_),
    .X(net506));
 sg13g2_buf_8 fanout507 (.A(_1864_),
    .X(net507));
 sg13g2_buf_8 fanout508 (.A(_1076_),
    .X(net508));
 sg13g2_buf_8 fanout509 (.A(_1043_),
    .X(net509));
 sg13g2_buf_8 fanout510 (.A(_0879_),
    .X(net510));
 sg13g2_buf_2 fanout511 (.A(_0879_),
    .X(net511));
 sg13g2_buf_8 fanout512 (.A(_0824_),
    .X(net512));
 sg13g2_buf_8 fanout513 (.A(_0813_),
    .X(net513));
 sg13g2_buf_8 fanout514 (.A(_0791_),
    .X(net514));
 sg13g2_buf_8 fanout515 (.A(_0780_),
    .X(net515));
 sg13g2_buf_8 fanout516 (.A(_0109_),
    .X(net516));
 sg13g2_buf_8 fanout517 (.A(_1955_),
    .X(net517));
 sg13g2_buf_2 fanout518 (.A(_1142_),
    .X(net518));
 sg13g2_buf_8 fanout519 (.A(net520),
    .X(net519));
 sg13g2_buf_8 fanout520 (.A(_0656_),
    .X(net520));
 sg13g2_buf_8 fanout521 (.A(_0655_),
    .X(net521));
 sg13g2_buf_8 fanout522 (.A(_2607_),
    .X(net522));
 sg13g2_buf_8 fanout523 (.A(net524),
    .X(net523));
 sg13g2_buf_8 fanout524 (.A(net525),
    .X(net524));
 sg13g2_buf_8 fanout525 (.A(_2588_),
    .X(net525));
 sg13g2_buf_8 fanout526 (.A(net528),
    .X(net526));
 sg13g2_buf_1 fanout527 (.A(net528),
    .X(net527));
 sg13g2_buf_8 fanout528 (.A(_2575_),
    .X(net528));
 sg13g2_buf_8 fanout529 (.A(net530),
    .X(net529));
 sg13g2_buf_8 fanout530 (.A(net531),
    .X(net530));
 sg13g2_buf_8 fanout531 (.A(_2574_),
    .X(net531));
 sg13g2_buf_8 fanout532 (.A(_1317_),
    .X(net532));
 sg13g2_buf_8 fanout533 (.A(_1229_),
    .X(net533));
 sg13g2_buf_8 fanout534 (.A(_1196_),
    .X(net534));
 sg13g2_buf_2 fanout535 (.A(_1196_),
    .X(net535));
 sg13g2_buf_8 fanout536 (.A(net537),
    .X(net536));
 sg13g2_buf_8 fanout537 (.A(_1185_),
    .X(net537));
 sg13g2_buf_8 fanout538 (.A(_1185_),
    .X(net538));
 sg13g2_buf_8 fanout539 (.A(_0560_),
    .X(net539));
 sg13g2_buf_8 fanout540 (.A(_1962_),
    .X(net540));
 sg13g2_buf_8 fanout541 (.A(_2603_),
    .X(net541));
 sg13g2_buf_8 fanout542 (.A(net543),
    .X(net542));
 sg13g2_buf_8 fanout543 (.A(_2589_),
    .X(net543));
 sg13g2_buf_8 fanout544 (.A(_2030_),
    .X(net544));
 sg13g2_buf_8 fanout545 (.A(_1306_),
    .X(net545));
 sg13g2_buf_8 fanout546 (.A(_1306_),
    .X(net546));
 sg13g2_buf_8 fanout547 (.A(_0934_),
    .X(net547));
 sg13g2_buf_8 fanout548 (.A(net549),
    .X(net548));
 sg13g2_buf_8 fanout549 (.A(_0571_),
    .X(net549));
 sg13g2_buf_8 fanout550 (.A(_0065_),
    .X(net550));
 sg13g2_buf_8 fanout551 (.A(_2745_),
    .X(net551));
 sg13g2_buf_8 fanout552 (.A(_2734_),
    .X(net552));
 sg13g2_buf_2 fanout553 (.A(_2734_),
    .X(net553));
 sg13g2_buf_8 fanout554 (.A(_2723_),
    .X(net554));
 sg13g2_buf_1 fanout555 (.A(_2723_),
    .X(net555));
 sg13g2_buf_8 fanout556 (.A(_2712_),
    .X(net556));
 sg13g2_buf_8 fanout557 (.A(_2701_),
    .X(net557));
 sg13g2_buf_8 fanout558 (.A(_2679_),
    .X(net558));
 sg13g2_buf_8 fanout559 (.A(_2646_),
    .X(net559));
 sg13g2_buf_8 fanout560 (.A(net561),
    .X(net560));
 sg13g2_buf_8 fanout561 (.A(_2602_),
    .X(net561));
 sg13g2_buf_8 fanout562 (.A(net564),
    .X(net562));
 sg13g2_buf_8 fanout563 (.A(net564),
    .X(net563));
 sg13g2_buf_8 fanout564 (.A(net565),
    .X(net564));
 sg13g2_buf_8 fanout565 (.A(_2558_),
    .X(net565));
 sg13g2_buf_8 fanout566 (.A(net569),
    .X(net566));
 sg13g2_buf_8 fanout567 (.A(net569),
    .X(net567));
 sg13g2_buf_8 fanout568 (.A(net569),
    .X(net568));
 sg13g2_buf_8 fanout569 (.A(net81),
    .X(net569));
 sg13g2_buf_8 fanout570 (.A(\flag.flag_abrosexual_inst.pix_y[8] ),
    .X(net570));
 sg13g2_buf_1 fanout571 (.A(\flag.flag_abrosexual_inst.pix_y[8] ),
    .X(net571));
 sg13g2_buf_8 fanout572 (.A(net574),
    .X(net572));
 sg13g2_buf_8 fanout573 (.A(net574),
    .X(net573));
 sg13g2_buf_2 fanout574 (.A(\flag.flag_abrosexual_inst.pix_y[7] ),
    .X(net574));
 sg13g2_buf_8 fanout575 (.A(net576),
    .X(net575));
 sg13g2_buf_8 fanout576 (.A(\flag.flag_abrosexual_inst.pix_y[7] ),
    .X(net576));
 sg13g2_buf_8 fanout577 (.A(net578),
    .X(net577));
 sg13g2_buf_8 fanout578 (.A(net579),
    .X(net578));
 sg13g2_buf_8 fanout579 (.A(net77),
    .X(net579));
 sg13g2_buf_8 fanout580 (.A(net581),
    .X(net580));
 sg13g2_buf_8 fanout581 (.A(\flag.flag_abrosexual_inst.pix_y[6] ),
    .X(net581));
 sg13g2_buf_8 fanout582 (.A(net584),
    .X(net582));
 sg13g2_buf_1 fanout583 (.A(net584),
    .X(net583));
 sg13g2_buf_8 fanout584 (.A(net75),
    .X(net584));
 sg13g2_buf_8 fanout585 (.A(net586),
    .X(net585));
 sg13g2_buf_8 fanout586 (.A(\flag.flag_abrosexual_inst.pix_y[5] ),
    .X(net586));
 sg13g2_buf_8 fanout587 (.A(net74),
    .X(net587));
 sg13g2_buf_1 fanout588 (.A(\flag.flag_abrosexual_inst.pix_y[4] ),
    .X(net588));
 sg13g2_buf_8 fanout589 (.A(net591),
    .X(net589));
 sg13g2_buf_2 fanout590 (.A(net591),
    .X(net590));
 sg13g2_buf_2 fanout591 (.A(\flag.flag_abrosexual_inst.pix_y[4] ),
    .X(net591));
 sg13g2_buf_8 fanout592 (.A(net593),
    .X(net592));
 sg13g2_buf_8 fanout593 (.A(net70),
    .X(net593));
 sg13g2_buf_2 fanout594 (.A(net70),
    .X(net594));
 sg13g2_buf_8 fanout595 (.A(net597),
    .X(net595));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596));
 sg13g2_buf_8 fanout597 (.A(net80),
    .X(net597));
 sg13g2_buf_8 fanout598 (.A(net78),
    .X(net598));
 sg13g2_buf_8 fanout599 (.A(\flag.flag_abrosexual_inst.pix_y[1] ),
    .X(net599));
 sg13g2_buf_8 fanout600 (.A(net605),
    .X(net600));
 sg13g2_buf_1 fanout601 (.A(net605),
    .X(net601));
 sg13g2_buf_8 fanout602 (.A(net605),
    .X(net602));
 sg13g2_buf_8 fanout603 (.A(net605),
    .X(net603));
 sg13g2_buf_1 fanout604 (.A(net605),
    .X(net604));
 sg13g2_buf_8 fanout605 (.A(\flag.flag_abrosexual_inst.pix_y[0] ),
    .X(net605));
 sg13g2_buf_8 fanout606 (.A(net609),
    .X(net606));
 sg13g2_buf_8 fanout607 (.A(net608),
    .X(net607));
 sg13g2_buf_8 fanout608 (.A(net609),
    .X(net608));
 sg13g2_buf_8 fanout609 (.A(net610),
    .X(net609));
 sg13g2_buf_2 fanout610 (.A(net73),
    .X(net610));
 sg13g2_buf_8 fanout611 (.A(net614),
    .X(net611));
 sg13g2_buf_8 fanout612 (.A(net613),
    .X(net612));
 sg13g2_buf_1 fanout613 (.A(net614),
    .X(net613));
 sg13g2_buf_8 fanout614 (.A(net615),
    .X(net614));
 sg13g2_buf_2 fanout615 (.A(net72),
    .X(net615));
 sg13g2_buf_8 fanout616 (.A(net619),
    .X(net616));
 sg13g2_buf_8 fanout617 (.A(net619),
    .X(net617));
 sg13g2_buf_8 fanout618 (.A(net619),
    .X(net618));
 sg13g2_buf_8 fanout619 (.A(net620),
    .X(net619));
 sg13g2_buf_8 fanout620 (.A(net67),
    .X(net620));
 sg13g2_buf_8 fanout621 (.A(net624),
    .X(net621));
 sg13g2_buf_8 fanout622 (.A(net624),
    .X(net622));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623));
 sg13g2_buf_8 fanout624 (.A(net625),
    .X(net624));
 sg13g2_buf_8 fanout625 (.A(net64),
    .X(net625));
 sg13g2_buf_8 fanout626 (.A(net630),
    .X(net626));
 sg13g2_buf_2 fanout627 (.A(net630),
    .X(net627));
 sg13g2_buf_8 fanout628 (.A(net630),
    .X(net628));
 sg13g2_buf_8 fanout629 (.A(net630),
    .X(net629));
 sg13g2_buf_8 fanout630 (.A(\flag.flag_abrosexual_inst.pix_x[5] ),
    .X(net630));
 sg13g2_buf_8 fanout631 (.A(net68),
    .X(net631));
 sg13g2_buf_8 fanout632 (.A(net635),
    .X(net632));
 sg13g2_buf_8 fanout633 (.A(net634),
    .X(net633));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634));
 sg13g2_buf_8 fanout635 (.A(net82),
    .X(net635));
 sg13g2_buf_8 fanout636 (.A(net638),
    .X(net636));
 sg13g2_buf_8 fanout637 (.A(net638),
    .X(net637));
 sg13g2_buf_8 fanout638 (.A(\flag.flag_abrosexual_inst.pix_x[3] ),
    .X(net638));
 sg13g2_buf_8 fanout639 (.A(net640),
    .X(net639));
 sg13g2_buf_8 fanout640 (.A(\flag.flag_abrosexual_inst.pix_x[2] ),
    .X(net640));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641));
 sg13g2_buf_8 fanout642 (.A(\flag.flag_abrosexual_inst.pix_x[2] ),
    .X(net642));
 sg13g2_buf_8 fanout643 (.A(net644),
    .X(net643));
 sg13g2_buf_1 fanout644 (.A(net645),
    .X(net644));
 sg13g2_buf_1 fanout645 (.A(\flag.flag_abrosexual_inst.pix_x[1] ),
    .X(net645));
 sg13g2_buf_8 fanout646 (.A(\flag.flag_abrosexual_inst.pix_x[1] ),
    .X(net646));
 sg13g2_buf_8 fanout647 (.A(net651),
    .X(net647));
 sg13g2_buf_8 fanout648 (.A(net650),
    .X(net648));
 sg13g2_buf_8 fanout649 (.A(net651),
    .X(net649));
 sg13g2_buf_2 fanout650 (.A(net651),
    .X(net650));
 sg13g2_buf_8 fanout651 (.A(net76),
    .X(net651));
 sg13g2_buf_8 fanout652 (.A(net653),
    .X(net652));
 sg13g2_buf_8 fanout653 (.A(\flag.flag_abrosexual_inst.pix_x[0] ),
    .X(net653));
 sg13g2_buf_8 fanout654 (.A(net655),
    .X(net654));
 sg13g2_buf_8 fanout655 (.A(net656),
    .X(net655));
 sg13g2_buf_8 fanout656 (.A(rst_n),
    .X(net656));
 sg13g2_buf_2 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[4]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[5]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[6]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[7]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(uio_in[0]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(uio_in[1]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(uio_in[2]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[3]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[4]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[5]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[6]),
    .X(net12));
 sg13g2_tielo tt_um_rebeccargb_vga_pride_13 (.L_LO(net13));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sg13g2_buf_1 clkload0 (.A(clknet_3_0__leaf_clk));
 sg13g2_buf_1 clkload1 (.A(clknet_3_1__leaf_clk));
 sg13g2_buf_1 clkload2 (.A(clknet_3_2__leaf_clk));
 sg13g2_buf_1 clkload3 (.A(clknet_3_3__leaf_clk));
 sg13g2_buf_1 clkload4 (.A(clknet_3_6__leaf_clk));
 sg13g2_buf_1 clkload5 (.A(clknet_3_7__leaf_clk));
 sg13g2_dlygate4sd3_1 hold1 (.A(\counter[3] ),
    .X(net51));
 sg13g2_dlygate4sd3_1 hold2 (.A(_0028_),
    .X(net52));
 sg13g2_dlygate4sd3_1 hold3 (.A(\counter[5] ),
    .X(net53));
 sg13g2_dlygate4sd3_1 hold4 (.A(_0030_),
    .X(net54));
 sg13g2_dlygate4sd3_1 hold5 (.A(\hvsync_gen.vpos[9] ),
    .X(net55));
 sg13g2_dlygate4sd3_1 hold6 (.A(\counter[6] ),
    .X(net56));
 sg13g2_dlygate4sd3_1 hold7 (.A(_2022_),
    .X(net57));
 sg13g2_dlygate4sd3_1 hold8 (.A(\counter[1] ),
    .X(net58));
 sg13g2_dlygate4sd3_1 hold9 (.A(_1987_),
    .X(net59));
 sg13g2_dlygate4sd3_1 hold10 (.A(\counter[2] ),
    .X(net60));
 sg13g2_dlygate4sd3_1 hold11 (.A(_0027_),
    .X(net61));
 sg13g2_dlygate4sd3_1 hold12 (.A(\counter[0] ),
    .X(net62));
 sg13g2_dlygate4sd3_1 hold13 (.A(_1973_),
    .X(net63));
 sg13g2_dlygate4sd3_1 hold14 (.A(\flag.flag_abrosexual_inst.pix_x[6] ),
    .X(net64));
 sg13g2_dlygate4sd3_1 hold15 (.A(\counter[4] ),
    .X(net65));
 sg13g2_dlygate4sd3_1 hold16 (.A(_0029_),
    .X(net66));
 sg13g2_dlygate4sd3_1 hold17 (.A(\flag.flag_abrosexual_inst.pix_x[7] ),
    .X(net67));
 sg13g2_dlygate4sd3_1 hold18 (.A(\flag.flag_abrosexual_inst.pix_x[5] ),
    .X(net68));
 sg13g2_dlygate4sd3_1 hold19 (.A(_1919_),
    .X(net69));
 sg13g2_dlygate4sd3_1 hold20 (.A(\flag.flag_abrosexual_inst.pix_y[3] ),
    .X(net70));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0014_),
    .X(net71));
 sg13g2_dlygate4sd3_1 hold22 (.A(\flag.flag_abrosexual_inst.pix_x[8] ),
    .X(net72));
 sg13g2_dlygate4sd3_1 hold23 (.A(\flag.flag_abrosexual_inst.pix_x[9] ),
    .X(net73));
 sg13g2_dlygate4sd3_1 hold24 (.A(\flag.flag_abrosexual_inst.pix_y[4] ),
    .X(net74));
 sg13g2_dlygate4sd3_1 hold25 (.A(\flag.flag_abrosexual_inst.pix_y[5] ),
    .X(net75));
 sg13g2_dlygate4sd3_1 hold26 (.A(\flag.flag_abrosexual_inst.pix_x[0] ),
    .X(net76));
 sg13g2_dlygate4sd3_1 hold27 (.A(\flag.flag_abrosexual_inst.pix_y[6] ),
    .X(net77));
 sg13g2_dlygate4sd3_1 hold28 (.A(\flag.flag_abrosexual_inst.pix_y[1] ),
    .X(net78));
 sg13g2_dlygate4sd3_1 hold29 (.A(_0016_),
    .X(net79));
 sg13g2_dlygate4sd3_1 hold30 (.A(\flag.flag_abrosexual_inst.pix_y[2] ),
    .X(net80));
 sg13g2_dlygate4sd3_1 hold31 (.A(\flag.flag_abrosexual_inst.pix_y[8] ),
    .X(net81));
 sg13g2_dlygate4sd3_1 hold32 (.A(\flag.flag_abrosexual_inst.pix_x[4] ),
    .X(net82));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_4 FILLER_0_238 ();
 sg13g2_fill_1 FILLER_0_242 ();
 sg13g2_decap_8 FILLER_0_251 ();
 sg13g2_decap_8 FILLER_0_258 ();
 sg13g2_fill_2 FILLER_0_265 ();
 sg13g2_fill_1 FILLER_0_271 ();
 sg13g2_decap_8 FILLER_0_276 ();
 sg13g2_decap_8 FILLER_0_283 ();
 sg13g2_decap_8 FILLER_0_290 ();
 sg13g2_decap_8 FILLER_0_297 ();
 sg13g2_decap_8 FILLER_0_304 ();
 sg13g2_decap_8 FILLER_0_311 ();
 sg13g2_decap_8 FILLER_0_318 ();
 sg13g2_decap_8 FILLER_0_325 ();
 sg13g2_decap_8 FILLER_0_332 ();
 sg13g2_decap_8 FILLER_0_339 ();
 sg13g2_decap_8 FILLER_0_346 ();
 sg13g2_decap_8 FILLER_0_353 ();
 sg13g2_decap_8 FILLER_0_360 ();
 sg13g2_decap_8 FILLER_0_367 ();
 sg13g2_decap_8 FILLER_0_374 ();
 sg13g2_decap_8 FILLER_0_381 ();
 sg13g2_decap_8 FILLER_0_388 ();
 sg13g2_decap_8 FILLER_0_395 ();
 sg13g2_decap_8 FILLER_0_402 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_4 FILLER_1_255 ();
 sg13g2_fill_2 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_282 ();
 sg13g2_decap_8 FILLER_1_289 ();
 sg13g2_decap_8 FILLER_1_296 ();
 sg13g2_decap_8 FILLER_1_303 ();
 sg13g2_decap_8 FILLER_1_310 ();
 sg13g2_decap_8 FILLER_1_317 ();
 sg13g2_decap_8 FILLER_1_324 ();
 sg13g2_decap_8 FILLER_1_331 ();
 sg13g2_decap_8 FILLER_1_338 ();
 sg13g2_decap_8 FILLER_1_345 ();
 sg13g2_decap_8 FILLER_1_352 ();
 sg13g2_decap_8 FILLER_1_359 ();
 sg13g2_decap_8 FILLER_1_366 ();
 sg13g2_decap_8 FILLER_1_373 ();
 sg13g2_decap_8 FILLER_1_380 ();
 sg13g2_decap_8 FILLER_1_387 ();
 sg13g2_decap_8 FILLER_1_394 ();
 sg13g2_decap_8 FILLER_1_401 ();
 sg13g2_fill_1 FILLER_1_408 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_8 FILLER_2_7 ();
 sg13g2_decap_8 FILLER_2_14 ();
 sg13g2_decap_8 FILLER_2_21 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_decap_8 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_63 ();
 sg13g2_decap_8 FILLER_2_70 ();
 sg13g2_decap_8 FILLER_2_77 ();
 sg13g2_decap_8 FILLER_2_84 ();
 sg13g2_decap_8 FILLER_2_91 ();
 sg13g2_decap_8 FILLER_2_98 ();
 sg13g2_decap_8 FILLER_2_105 ();
 sg13g2_decap_8 FILLER_2_112 ();
 sg13g2_decap_8 FILLER_2_119 ();
 sg13g2_decap_8 FILLER_2_126 ();
 sg13g2_decap_8 FILLER_2_133 ();
 sg13g2_decap_8 FILLER_2_140 ();
 sg13g2_decap_8 FILLER_2_147 ();
 sg13g2_decap_8 FILLER_2_154 ();
 sg13g2_decap_8 FILLER_2_161 ();
 sg13g2_decap_8 FILLER_2_168 ();
 sg13g2_decap_8 FILLER_2_175 ();
 sg13g2_decap_8 FILLER_2_182 ();
 sg13g2_decap_8 FILLER_2_189 ();
 sg13g2_decap_8 FILLER_2_196 ();
 sg13g2_decap_4 FILLER_2_203 ();
 sg13g2_fill_1 FILLER_2_207 ();
 sg13g2_fill_1 FILLER_2_238 ();
 sg13g2_fill_2 FILLER_2_247 ();
 sg13g2_fill_1 FILLER_2_249 ();
 sg13g2_fill_2 FILLER_2_279 ();
 sg13g2_fill_1 FILLER_2_281 ();
 sg13g2_decap_8 FILLER_2_297 ();
 sg13g2_decap_8 FILLER_2_304 ();
 sg13g2_decap_8 FILLER_2_311 ();
 sg13g2_decap_8 FILLER_2_318 ();
 sg13g2_decap_8 FILLER_2_325 ();
 sg13g2_decap_8 FILLER_2_332 ();
 sg13g2_decap_8 FILLER_2_339 ();
 sg13g2_decap_8 FILLER_2_346 ();
 sg13g2_decap_8 FILLER_2_353 ();
 sg13g2_decap_8 FILLER_2_360 ();
 sg13g2_decap_8 FILLER_2_367 ();
 sg13g2_decap_8 FILLER_2_374 ();
 sg13g2_decap_8 FILLER_2_381 ();
 sg13g2_decap_8 FILLER_2_388 ();
 sg13g2_decap_8 FILLER_2_395 ();
 sg13g2_decap_8 FILLER_2_402 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_fill_2 FILLER_3_196 ();
 sg13g2_fill_1 FILLER_3_198 ();
 sg13g2_fill_1 FILLER_3_224 ();
 sg13g2_fill_2 FILLER_3_241 ();
 sg13g2_fill_1 FILLER_3_243 ();
 sg13g2_decap_8 FILLER_3_249 ();
 sg13g2_decap_4 FILLER_3_256 ();
 sg13g2_fill_2 FILLER_3_291 ();
 sg13g2_fill_1 FILLER_3_293 ();
 sg13g2_decap_8 FILLER_3_304 ();
 sg13g2_decap_8 FILLER_3_311 ();
 sg13g2_decap_8 FILLER_3_318 ();
 sg13g2_decap_8 FILLER_3_325 ();
 sg13g2_decap_8 FILLER_3_332 ();
 sg13g2_decap_8 FILLER_3_339 ();
 sg13g2_decap_8 FILLER_3_346 ();
 sg13g2_decap_8 FILLER_3_353 ();
 sg13g2_decap_8 FILLER_3_360 ();
 sg13g2_decap_8 FILLER_3_367 ();
 sg13g2_decap_8 FILLER_3_374 ();
 sg13g2_decap_8 FILLER_3_381 ();
 sg13g2_decap_8 FILLER_3_388 ();
 sg13g2_decap_8 FILLER_3_395 ();
 sg13g2_decap_8 FILLER_3_402 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_fill_2 FILLER_4_196 ();
 sg13g2_fill_2 FILLER_4_214 ();
 sg13g2_fill_1 FILLER_4_216 ();
 sg13g2_decap_8 FILLER_4_253 ();
 sg13g2_decap_4 FILLER_4_260 ();
 sg13g2_fill_1 FILLER_4_269 ();
 sg13g2_decap_4 FILLER_4_274 ();
 sg13g2_decap_8 FILLER_4_303 ();
 sg13g2_decap_8 FILLER_4_310 ();
 sg13g2_decap_8 FILLER_4_317 ();
 sg13g2_decap_8 FILLER_4_324 ();
 sg13g2_decap_8 FILLER_4_331 ();
 sg13g2_decap_8 FILLER_4_338 ();
 sg13g2_decap_8 FILLER_4_345 ();
 sg13g2_decap_8 FILLER_4_352 ();
 sg13g2_decap_8 FILLER_4_359 ();
 sg13g2_decap_8 FILLER_4_366 ();
 sg13g2_decap_8 FILLER_4_373 ();
 sg13g2_decap_8 FILLER_4_380 ();
 sg13g2_decap_8 FILLER_4_387 ();
 sg13g2_decap_8 FILLER_4_394 ();
 sg13g2_decap_8 FILLER_4_401 ();
 sg13g2_fill_1 FILLER_4_408 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_7 ();
 sg13g2_decap_8 FILLER_5_14 ();
 sg13g2_decap_8 FILLER_5_21 ();
 sg13g2_decap_8 FILLER_5_28 ();
 sg13g2_decap_8 FILLER_5_35 ();
 sg13g2_decap_8 FILLER_5_42 ();
 sg13g2_decap_8 FILLER_5_49 ();
 sg13g2_decap_8 FILLER_5_56 ();
 sg13g2_decap_8 FILLER_5_63 ();
 sg13g2_decap_8 FILLER_5_70 ();
 sg13g2_decap_8 FILLER_5_77 ();
 sg13g2_decap_8 FILLER_5_84 ();
 sg13g2_decap_8 FILLER_5_91 ();
 sg13g2_decap_8 FILLER_5_98 ();
 sg13g2_decap_8 FILLER_5_105 ();
 sg13g2_decap_8 FILLER_5_112 ();
 sg13g2_decap_8 FILLER_5_119 ();
 sg13g2_decap_8 FILLER_5_126 ();
 sg13g2_decap_8 FILLER_5_133 ();
 sg13g2_decap_8 FILLER_5_140 ();
 sg13g2_decap_8 FILLER_5_147 ();
 sg13g2_decap_8 FILLER_5_154 ();
 sg13g2_decap_8 FILLER_5_161 ();
 sg13g2_decap_8 FILLER_5_168 ();
 sg13g2_decap_8 FILLER_5_175 ();
 sg13g2_decap_8 FILLER_5_182 ();
 sg13g2_decap_8 FILLER_5_189 ();
 sg13g2_fill_1 FILLER_5_222 ();
 sg13g2_decap_8 FILLER_5_248 ();
 sg13g2_decap_4 FILLER_5_255 ();
 sg13g2_fill_1 FILLER_5_259 ();
 sg13g2_fill_1 FILLER_5_278 ();
 sg13g2_decap_8 FILLER_5_304 ();
 sg13g2_decap_8 FILLER_5_311 ();
 sg13g2_decap_8 FILLER_5_318 ();
 sg13g2_decap_8 FILLER_5_325 ();
 sg13g2_decap_8 FILLER_5_332 ();
 sg13g2_decap_8 FILLER_5_339 ();
 sg13g2_decap_8 FILLER_5_346 ();
 sg13g2_decap_8 FILLER_5_353 ();
 sg13g2_decap_8 FILLER_5_360 ();
 sg13g2_decap_8 FILLER_5_367 ();
 sg13g2_decap_8 FILLER_5_374 ();
 sg13g2_decap_8 FILLER_5_381 ();
 sg13g2_decap_8 FILLER_5_388 ();
 sg13g2_decap_8 FILLER_5_395 ();
 sg13g2_decap_8 FILLER_5_402 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_fill_2 FILLER_6_154 ();
 sg13g2_fill_1 FILLER_6_156 ();
 sg13g2_decap_8 FILLER_6_211 ();
 sg13g2_decap_8 FILLER_6_222 ();
 sg13g2_decap_8 FILLER_6_229 ();
 sg13g2_fill_2 FILLER_6_236 ();
 sg13g2_fill_2 FILLER_6_248 ();
 sg13g2_fill_2 FILLER_6_258 ();
 sg13g2_decap_4 FILLER_6_280 ();
 sg13g2_fill_2 FILLER_6_284 ();
 sg13g2_decap_8 FILLER_6_295 ();
 sg13g2_decap_8 FILLER_6_302 ();
 sg13g2_decap_8 FILLER_6_309 ();
 sg13g2_decap_8 FILLER_6_316 ();
 sg13g2_decap_8 FILLER_6_323 ();
 sg13g2_decap_8 FILLER_6_330 ();
 sg13g2_decap_8 FILLER_6_337 ();
 sg13g2_decap_8 FILLER_6_344 ();
 sg13g2_decap_8 FILLER_6_351 ();
 sg13g2_decap_8 FILLER_6_358 ();
 sg13g2_decap_8 FILLER_6_365 ();
 sg13g2_decap_8 FILLER_6_372 ();
 sg13g2_decap_8 FILLER_6_379 ();
 sg13g2_decap_8 FILLER_6_386 ();
 sg13g2_decap_8 FILLER_6_393 ();
 sg13g2_decap_8 FILLER_6_400 ();
 sg13g2_fill_2 FILLER_6_407 ();
 sg13g2_decap_8 FILLER_7_0 ();
 sg13g2_decap_8 FILLER_7_7 ();
 sg13g2_decap_8 FILLER_7_14 ();
 sg13g2_decap_8 FILLER_7_21 ();
 sg13g2_decap_8 FILLER_7_28 ();
 sg13g2_decap_8 FILLER_7_35 ();
 sg13g2_decap_8 FILLER_7_42 ();
 sg13g2_decap_8 FILLER_7_49 ();
 sg13g2_decap_8 FILLER_7_56 ();
 sg13g2_decap_8 FILLER_7_63 ();
 sg13g2_decap_8 FILLER_7_70 ();
 sg13g2_decap_8 FILLER_7_77 ();
 sg13g2_decap_8 FILLER_7_84 ();
 sg13g2_decap_8 FILLER_7_91 ();
 sg13g2_decap_8 FILLER_7_98 ();
 sg13g2_decap_8 FILLER_7_105 ();
 sg13g2_decap_8 FILLER_7_112 ();
 sg13g2_decap_8 FILLER_7_119 ();
 sg13g2_decap_8 FILLER_7_126 ();
 sg13g2_fill_2 FILLER_7_133 ();
 sg13g2_fill_1 FILLER_7_135 ();
 sg13g2_decap_8 FILLER_7_140 ();
 sg13g2_decap_8 FILLER_7_147 ();
 sg13g2_fill_2 FILLER_7_163 ();
 sg13g2_fill_2 FILLER_7_201 ();
 sg13g2_fill_1 FILLER_7_203 ();
 sg13g2_decap_8 FILLER_7_208 ();
 sg13g2_decap_4 FILLER_7_215 ();
 sg13g2_fill_1 FILLER_7_219 ();
 sg13g2_fill_2 FILLER_7_228 ();
 sg13g2_fill_2 FILLER_7_258 ();
 sg13g2_fill_1 FILLER_7_260 ();
 sg13g2_decap_8 FILLER_7_271 ();
 sg13g2_decap_8 FILLER_7_278 ();
 sg13g2_decap_8 FILLER_7_285 ();
 sg13g2_decap_8 FILLER_7_292 ();
 sg13g2_decap_8 FILLER_7_299 ();
 sg13g2_decap_8 FILLER_7_306 ();
 sg13g2_decap_8 FILLER_7_313 ();
 sg13g2_decap_8 FILLER_7_320 ();
 sg13g2_decap_8 FILLER_7_327 ();
 sg13g2_decap_8 FILLER_7_334 ();
 sg13g2_decap_8 FILLER_7_341 ();
 sg13g2_decap_8 FILLER_7_348 ();
 sg13g2_decap_8 FILLER_7_355 ();
 sg13g2_decap_8 FILLER_7_362 ();
 sg13g2_decap_8 FILLER_7_369 ();
 sg13g2_decap_8 FILLER_7_376 ();
 sg13g2_decap_8 FILLER_7_383 ();
 sg13g2_decap_8 FILLER_7_390 ();
 sg13g2_decap_8 FILLER_7_397 ();
 sg13g2_decap_4 FILLER_7_404 ();
 sg13g2_fill_1 FILLER_7_408 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_4 FILLER_8_126 ();
 sg13g2_fill_1 FILLER_8_174 ();
 sg13g2_fill_1 FILLER_8_180 ();
 sg13g2_fill_1 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_242 ();
 sg13g2_fill_2 FILLER_8_249 ();
 sg13g2_fill_1 FILLER_8_251 ();
 sg13g2_fill_1 FILLER_8_285 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_fill_2 FILLER_8_406 ();
 sg13g2_fill_1 FILLER_8_408 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_fill_2 FILLER_9_133 ();
 sg13g2_fill_1 FILLER_9_135 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_178 ();
 sg13g2_fill_1 FILLER_9_189 ();
 sg13g2_fill_2 FILLER_9_203 ();
 sg13g2_fill_2 FILLER_9_234 ();
 sg13g2_decap_8 FILLER_9_255 ();
 sg13g2_decap_4 FILLER_9_262 ();
 sg13g2_fill_1 FILLER_9_269 ();
 sg13g2_decap_8 FILLER_9_300 ();
 sg13g2_decap_8 FILLER_9_307 ();
 sg13g2_decap_8 FILLER_9_314 ();
 sg13g2_decap_8 FILLER_9_321 ();
 sg13g2_decap_8 FILLER_9_328 ();
 sg13g2_decap_8 FILLER_9_335 ();
 sg13g2_decap_8 FILLER_9_342 ();
 sg13g2_decap_8 FILLER_9_349 ();
 sg13g2_decap_8 FILLER_9_356 ();
 sg13g2_decap_8 FILLER_9_363 ();
 sg13g2_decap_8 FILLER_9_370 ();
 sg13g2_decap_8 FILLER_9_377 ();
 sg13g2_decap_8 FILLER_9_384 ();
 sg13g2_decap_8 FILLER_9_391 ();
 sg13g2_decap_8 FILLER_9_398 ();
 sg13g2_decap_4 FILLER_9_405 ();
 sg13g2_decap_8 FILLER_10_0 ();
 sg13g2_decap_8 FILLER_10_7 ();
 sg13g2_decap_8 FILLER_10_14 ();
 sg13g2_decap_8 FILLER_10_21 ();
 sg13g2_decap_8 FILLER_10_28 ();
 sg13g2_decap_8 FILLER_10_35 ();
 sg13g2_fill_1 FILLER_10_42 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_fill_1 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_58 ();
 sg13g2_fill_1 FILLER_10_78 ();
 sg13g2_decap_8 FILLER_10_89 ();
 sg13g2_decap_8 FILLER_10_96 ();
 sg13g2_decap_8 FILLER_10_103 ();
 sg13g2_decap_8 FILLER_10_110 ();
 sg13g2_decap_8 FILLER_10_117 ();
 sg13g2_decap_8 FILLER_10_124 ();
 sg13g2_decap_8 FILLER_10_131 ();
 sg13g2_decap_4 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_142 ();
 sg13g2_fill_1 FILLER_10_184 ();
 sg13g2_decap_4 FILLER_10_194 ();
 sg13g2_fill_1 FILLER_10_198 ();
 sg13g2_fill_2 FILLER_10_219 ();
 sg13g2_decap_4 FILLER_10_240 ();
 sg13g2_fill_1 FILLER_10_282 ();
 sg13g2_decap_8 FILLER_10_304 ();
 sg13g2_decap_8 FILLER_10_311 ();
 sg13g2_decap_8 FILLER_10_318 ();
 sg13g2_decap_8 FILLER_10_325 ();
 sg13g2_decap_8 FILLER_10_332 ();
 sg13g2_decap_8 FILLER_10_339 ();
 sg13g2_decap_8 FILLER_10_346 ();
 sg13g2_decap_8 FILLER_10_353 ();
 sg13g2_decap_8 FILLER_10_360 ();
 sg13g2_decap_8 FILLER_10_367 ();
 sg13g2_decap_8 FILLER_10_374 ();
 sg13g2_decap_8 FILLER_10_381 ();
 sg13g2_decap_8 FILLER_10_388 ();
 sg13g2_decap_8 FILLER_10_395 ();
 sg13g2_decap_8 FILLER_10_402 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_fill_2 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_94 ();
 sg13g2_decap_8 FILLER_11_101 ();
 sg13g2_decap_8 FILLER_11_108 ();
 sg13g2_decap_8 FILLER_11_115 ();
 sg13g2_decap_8 FILLER_11_122 ();
 sg13g2_decap_4 FILLER_11_129 ();
 sg13g2_fill_2 FILLER_11_133 ();
 sg13g2_fill_1 FILLER_11_167 ();
 sg13g2_fill_2 FILLER_11_175 ();
 sg13g2_fill_2 FILLER_11_190 ();
 sg13g2_decap_4 FILLER_11_205 ();
 sg13g2_fill_2 FILLER_11_209 ();
 sg13g2_decap_4 FILLER_11_216 ();
 sg13g2_fill_1 FILLER_11_220 ();
 sg13g2_decap_8 FILLER_11_226 ();
 sg13g2_decap_4 FILLER_11_233 ();
 sg13g2_decap_8 FILLER_11_243 ();
 sg13g2_fill_1 FILLER_11_250 ();
 sg13g2_fill_1 FILLER_11_279 ();
 sg13g2_decap_4 FILLER_11_288 ();
 sg13g2_fill_1 FILLER_11_292 ();
 sg13g2_decap_8 FILLER_11_298 ();
 sg13g2_decap_8 FILLER_11_305 ();
 sg13g2_decap_8 FILLER_11_312 ();
 sg13g2_decap_8 FILLER_11_319 ();
 sg13g2_decap_8 FILLER_11_326 ();
 sg13g2_decap_8 FILLER_11_333 ();
 sg13g2_decap_8 FILLER_11_340 ();
 sg13g2_decap_8 FILLER_11_347 ();
 sg13g2_decap_8 FILLER_11_354 ();
 sg13g2_decap_8 FILLER_11_361 ();
 sg13g2_decap_8 FILLER_11_368 ();
 sg13g2_decap_8 FILLER_11_375 ();
 sg13g2_decap_8 FILLER_11_382 ();
 sg13g2_decap_8 FILLER_11_389 ();
 sg13g2_decap_8 FILLER_11_396 ();
 sg13g2_decap_4 FILLER_11_403 ();
 sg13g2_fill_2 FILLER_11_407 ();
 sg13g2_decap_8 FILLER_12_0 ();
 sg13g2_decap_8 FILLER_12_7 ();
 sg13g2_decap_8 FILLER_12_14 ();
 sg13g2_decap_8 FILLER_12_21 ();
 sg13g2_fill_2 FILLER_12_28 ();
 sg13g2_fill_1 FILLER_12_30 ();
 sg13g2_fill_2 FILLER_12_50 ();
 sg13g2_fill_2 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_106 ();
 sg13g2_decap_8 FILLER_12_113 ();
 sg13g2_decap_8 FILLER_12_120 ();
 sg13g2_fill_2 FILLER_12_127 ();
 sg13g2_fill_1 FILLER_12_129 ();
 sg13g2_fill_1 FILLER_12_179 ();
 sg13g2_fill_2 FILLER_12_216 ();
 sg13g2_fill_2 FILLER_12_235 ();
 sg13g2_fill_1 FILLER_12_237 ();
 sg13g2_fill_1 FILLER_12_251 ();
 sg13g2_fill_1 FILLER_12_260 ();
 sg13g2_decap_8 FILLER_12_294 ();
 sg13g2_decap_8 FILLER_12_301 ();
 sg13g2_decap_8 FILLER_12_308 ();
 sg13g2_decap_8 FILLER_12_315 ();
 sg13g2_decap_8 FILLER_12_322 ();
 sg13g2_decap_8 FILLER_12_329 ();
 sg13g2_decap_8 FILLER_12_336 ();
 sg13g2_decap_8 FILLER_12_343 ();
 sg13g2_decap_8 FILLER_12_350 ();
 sg13g2_decap_8 FILLER_12_357 ();
 sg13g2_decap_8 FILLER_12_364 ();
 sg13g2_decap_8 FILLER_12_371 ();
 sg13g2_decap_8 FILLER_12_378 ();
 sg13g2_decap_8 FILLER_12_385 ();
 sg13g2_decap_8 FILLER_12_392 ();
 sg13g2_decap_8 FILLER_12_399 ();
 sg13g2_fill_2 FILLER_12_406 ();
 sg13g2_fill_1 FILLER_12_408 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_fill_2 FILLER_13_35 ();
 sg13g2_fill_1 FILLER_13_37 ();
 sg13g2_fill_2 FILLER_13_61 ();
 sg13g2_fill_2 FILLER_13_81 ();
 sg13g2_decap_8 FILLER_13_113 ();
 sg13g2_fill_1 FILLER_13_124 ();
 sg13g2_fill_2 FILLER_13_227 ();
 sg13g2_fill_1 FILLER_13_229 ();
 sg13g2_fill_2 FILLER_13_260 ();
 sg13g2_fill_1 FILLER_13_267 ();
 sg13g2_fill_2 FILLER_13_276 ();
 sg13g2_fill_1 FILLER_13_278 ();
 sg13g2_fill_2 FILLER_13_287 ();
 sg13g2_fill_1 FILLER_13_289 ();
 sg13g2_decap_8 FILLER_13_298 ();
 sg13g2_decap_8 FILLER_13_305 ();
 sg13g2_decap_8 FILLER_13_312 ();
 sg13g2_decap_8 FILLER_13_319 ();
 sg13g2_decap_8 FILLER_13_326 ();
 sg13g2_decap_8 FILLER_13_333 ();
 sg13g2_decap_8 FILLER_13_340 ();
 sg13g2_decap_8 FILLER_13_347 ();
 sg13g2_decap_8 FILLER_13_354 ();
 sg13g2_decap_8 FILLER_13_361 ();
 sg13g2_decap_8 FILLER_13_368 ();
 sg13g2_decap_8 FILLER_13_375 ();
 sg13g2_decap_8 FILLER_13_382 ();
 sg13g2_decap_8 FILLER_13_389 ();
 sg13g2_decap_8 FILLER_13_396 ();
 sg13g2_decap_4 FILLER_13_403 ();
 sg13g2_fill_2 FILLER_13_407 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_4 FILLER_14_28 ();
 sg13g2_fill_1 FILLER_14_32 ();
 sg13g2_fill_2 FILLER_14_46 ();
 sg13g2_decap_4 FILLER_14_52 ();
 sg13g2_fill_2 FILLER_14_76 ();
 sg13g2_fill_1 FILLER_14_78 ();
 sg13g2_decap_4 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_fill_2 FILLER_14_112 ();
 sg13g2_fill_1 FILLER_14_114 ();
 sg13g2_fill_1 FILLER_14_162 ();
 sg13g2_decap_4 FILLER_14_202 ();
 sg13g2_fill_1 FILLER_14_210 ();
 sg13g2_fill_1 FILLER_14_224 ();
 sg13g2_fill_2 FILLER_14_246 ();
 sg13g2_fill_1 FILLER_14_256 ();
 sg13g2_decap_8 FILLER_14_292 ();
 sg13g2_decap_8 FILLER_14_299 ();
 sg13g2_decap_8 FILLER_14_306 ();
 sg13g2_decap_8 FILLER_14_313 ();
 sg13g2_decap_8 FILLER_14_320 ();
 sg13g2_decap_8 FILLER_14_327 ();
 sg13g2_decap_8 FILLER_14_334 ();
 sg13g2_decap_8 FILLER_14_341 ();
 sg13g2_decap_8 FILLER_14_348 ();
 sg13g2_decap_8 FILLER_14_355 ();
 sg13g2_decap_8 FILLER_14_362 ();
 sg13g2_decap_8 FILLER_14_369 ();
 sg13g2_decap_8 FILLER_14_376 ();
 sg13g2_decap_8 FILLER_14_383 ();
 sg13g2_decap_8 FILLER_14_390 ();
 sg13g2_decap_8 FILLER_14_397 ();
 sg13g2_decap_4 FILLER_14_404 ();
 sg13g2_fill_1 FILLER_14_408 ();
 sg13g2_decap_8 FILLER_15_0 ();
 sg13g2_decap_8 FILLER_15_7 ();
 sg13g2_decap_8 FILLER_15_14 ();
 sg13g2_decap_4 FILLER_15_21 ();
 sg13g2_fill_2 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_4 FILLER_15_60 ();
 sg13g2_decap_4 FILLER_15_69 ();
 sg13g2_fill_1 FILLER_15_73 ();
 sg13g2_fill_2 FILLER_15_90 ();
 sg13g2_fill_1 FILLER_15_92 ();
 sg13g2_decap_8 FILLER_15_105 ();
 sg13g2_decap_8 FILLER_15_112 ();
 sg13g2_decap_8 FILLER_15_119 ();
 sg13g2_decap_4 FILLER_15_126 ();
 sg13g2_fill_2 FILLER_15_130 ();
 sg13g2_decap_4 FILLER_15_159 ();
 sg13g2_fill_1 FILLER_15_163 ();
 sg13g2_decap_8 FILLER_15_217 ();
 sg13g2_fill_2 FILLER_15_228 ();
 sg13g2_fill_1 FILLER_15_230 ();
 sg13g2_fill_2 FILLER_15_244 ();
 sg13g2_fill_1 FILLER_15_246 ();
 sg13g2_fill_2 FILLER_15_252 ();
 sg13g2_fill_2 FILLER_15_258 ();
 sg13g2_decap_8 FILLER_15_265 ();
 sg13g2_decap_8 FILLER_15_272 ();
 sg13g2_fill_2 FILLER_15_279 ();
 sg13g2_fill_1 FILLER_15_281 ();
 sg13g2_decap_4 FILLER_15_290 ();
 sg13g2_fill_2 FILLER_15_294 ();
 sg13g2_decap_8 FILLER_15_299 ();
 sg13g2_decap_8 FILLER_15_306 ();
 sg13g2_decap_8 FILLER_15_313 ();
 sg13g2_decap_8 FILLER_15_320 ();
 sg13g2_decap_8 FILLER_15_327 ();
 sg13g2_decap_8 FILLER_15_334 ();
 sg13g2_decap_8 FILLER_15_341 ();
 sg13g2_decap_8 FILLER_15_348 ();
 sg13g2_decap_8 FILLER_15_355 ();
 sg13g2_decap_8 FILLER_15_362 ();
 sg13g2_decap_8 FILLER_15_369 ();
 sg13g2_decap_8 FILLER_15_376 ();
 sg13g2_decap_8 FILLER_15_383 ();
 sg13g2_decap_8 FILLER_15_390 ();
 sg13g2_decap_8 FILLER_15_397 ();
 sg13g2_decap_4 FILLER_15_404 ();
 sg13g2_fill_1 FILLER_15_408 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_fill_2 FILLER_16_28 ();
 sg13g2_fill_1 FILLER_16_30 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_4 FILLER_16_63 ();
 sg13g2_fill_1 FILLER_16_67 ();
 sg13g2_decap_4 FILLER_16_94 ();
 sg13g2_decap_8 FILLER_16_103 ();
 sg13g2_fill_2 FILLER_16_110 ();
 sg13g2_fill_1 FILLER_16_112 ();
 sg13g2_decap_4 FILLER_16_141 ();
 sg13g2_fill_1 FILLER_16_156 ();
 sg13g2_fill_2 FILLER_16_192 ();
 sg13g2_fill_1 FILLER_16_194 ();
 sg13g2_decap_8 FILLER_16_248 ();
 sg13g2_fill_2 FILLER_16_259 ();
 sg13g2_decap_4 FILLER_16_275 ();
 sg13g2_fill_2 FILLER_16_279 ();
 sg13g2_fill_1 FILLER_16_286 ();
 sg13g2_decap_8 FILLER_16_295 ();
 sg13g2_decap_8 FILLER_16_302 ();
 sg13g2_decap_8 FILLER_16_309 ();
 sg13g2_decap_8 FILLER_16_316 ();
 sg13g2_decap_8 FILLER_16_323 ();
 sg13g2_decap_8 FILLER_16_330 ();
 sg13g2_decap_8 FILLER_16_337 ();
 sg13g2_decap_8 FILLER_16_344 ();
 sg13g2_decap_8 FILLER_16_351 ();
 sg13g2_decap_8 FILLER_16_358 ();
 sg13g2_decap_8 FILLER_16_365 ();
 sg13g2_decap_8 FILLER_16_372 ();
 sg13g2_decap_8 FILLER_16_379 ();
 sg13g2_decap_8 FILLER_16_386 ();
 sg13g2_decap_8 FILLER_16_393 ();
 sg13g2_decap_8 FILLER_16_400 ();
 sg13g2_fill_2 FILLER_16_407 ();
 sg13g2_decap_8 FILLER_17_0 ();
 sg13g2_decap_8 FILLER_17_7 ();
 sg13g2_decap_8 FILLER_17_14 ();
 sg13g2_decap_8 FILLER_17_21 ();
 sg13g2_decap_8 FILLER_17_28 ();
 sg13g2_decap_4 FILLER_17_35 ();
 sg13g2_fill_2 FILLER_17_39 ();
 sg13g2_fill_2 FILLER_17_53 ();
 sg13g2_fill_1 FILLER_17_55 ();
 sg13g2_decap_4 FILLER_17_69 ();
 sg13g2_decap_4 FILLER_17_86 ();
 sg13g2_decap_8 FILLER_17_111 ();
 sg13g2_fill_2 FILLER_17_122 ();
 sg13g2_fill_1 FILLER_17_124 ();
 sg13g2_fill_1 FILLER_17_156 ();
 sg13g2_fill_2 FILLER_17_194 ();
 sg13g2_fill_1 FILLER_17_196 ();
 sg13g2_decap_4 FILLER_17_238 ();
 sg13g2_fill_2 FILLER_17_246 ();
 sg13g2_fill_1 FILLER_17_248 ();
 sg13g2_decap_4 FILLER_17_278 ();
 sg13g2_decap_8 FILLER_17_300 ();
 sg13g2_decap_8 FILLER_17_307 ();
 sg13g2_decap_8 FILLER_17_314 ();
 sg13g2_decap_8 FILLER_17_321 ();
 sg13g2_decap_8 FILLER_17_328 ();
 sg13g2_decap_8 FILLER_17_335 ();
 sg13g2_decap_8 FILLER_17_342 ();
 sg13g2_decap_8 FILLER_17_349 ();
 sg13g2_decap_8 FILLER_17_356 ();
 sg13g2_decap_8 FILLER_17_363 ();
 sg13g2_decap_8 FILLER_17_370 ();
 sg13g2_decap_8 FILLER_17_377 ();
 sg13g2_decap_8 FILLER_17_384 ();
 sg13g2_decap_8 FILLER_17_391 ();
 sg13g2_decap_8 FILLER_17_398 ();
 sg13g2_decap_4 FILLER_17_405 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_4 FILLER_18_21 ();
 sg13g2_fill_1 FILLER_18_25 ();
 sg13g2_decap_4 FILLER_18_34 ();
 sg13g2_fill_1 FILLER_18_38 ();
 sg13g2_decap_8 FILLER_18_47 ();
 sg13g2_fill_2 FILLER_18_81 ();
 sg13g2_fill_1 FILLER_18_108 ();
 sg13g2_fill_2 FILLER_18_141 ();
 sg13g2_fill_1 FILLER_18_151 ();
 sg13g2_decap_4 FILLER_18_176 ();
 sg13g2_decap_4 FILLER_18_186 ();
 sg13g2_fill_2 FILLER_18_206 ();
 sg13g2_fill_2 FILLER_18_230 ();
 sg13g2_fill_1 FILLER_18_245 ();
 sg13g2_fill_1 FILLER_18_267 ();
 sg13g2_fill_2 FILLER_18_281 ();
 sg13g2_decap_8 FILLER_18_300 ();
 sg13g2_decap_8 FILLER_18_307 ();
 sg13g2_decap_8 FILLER_18_314 ();
 sg13g2_decap_8 FILLER_18_321 ();
 sg13g2_decap_8 FILLER_18_328 ();
 sg13g2_fill_1 FILLER_18_335 ();
 sg13g2_fill_1 FILLER_18_340 ();
 sg13g2_decap_8 FILLER_18_345 ();
 sg13g2_decap_8 FILLER_18_352 ();
 sg13g2_decap_8 FILLER_18_359 ();
 sg13g2_decap_8 FILLER_18_366 ();
 sg13g2_decap_8 FILLER_18_373 ();
 sg13g2_decap_8 FILLER_18_380 ();
 sg13g2_decap_8 FILLER_18_387 ();
 sg13g2_decap_8 FILLER_18_394 ();
 sg13g2_decap_8 FILLER_18_401 ();
 sg13g2_fill_1 FILLER_18_408 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_4 FILLER_19_14 ();
 sg13g2_fill_2 FILLER_19_31 ();
 sg13g2_fill_1 FILLER_19_33 ();
 sg13g2_fill_2 FILLER_19_47 ();
 sg13g2_decap_4 FILLER_19_78 ();
 sg13g2_fill_2 FILLER_19_90 ();
 sg13g2_fill_1 FILLER_19_92 ();
 sg13g2_decap_4 FILLER_19_101 ();
 sg13g2_fill_2 FILLER_19_152 ();
 sg13g2_fill_1 FILLER_19_154 ();
 sg13g2_fill_1 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_221 ();
 sg13g2_fill_1 FILLER_19_228 ();
 sg13g2_decap_8 FILLER_19_288 ();
 sg13g2_decap_8 FILLER_19_295 ();
 sg13g2_decap_4 FILLER_19_302 ();
 sg13g2_fill_1 FILLER_19_306 ();
 sg13g2_decap_4 FILLER_19_321 ();
 sg13g2_fill_2 FILLER_19_325 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_fill_2 FILLER_19_406 ();
 sg13g2_fill_1 FILLER_19_408 ();
 sg13g2_decap_8 FILLER_20_0 ();
 sg13g2_decap_4 FILLER_20_7 ();
 sg13g2_decap_8 FILLER_20_48 ();
 sg13g2_decap_8 FILLER_20_55 ();
 sg13g2_decap_8 FILLER_20_62 ();
 sg13g2_decap_4 FILLER_20_69 ();
 sg13g2_fill_2 FILLER_20_73 ();
 sg13g2_decap_8 FILLER_20_96 ();
 sg13g2_decap_8 FILLER_20_103 ();
 sg13g2_fill_2 FILLER_20_110 ();
 sg13g2_fill_1 FILLER_20_112 ();
 sg13g2_decap_8 FILLER_20_119 ();
 sg13g2_fill_2 FILLER_20_126 ();
 sg13g2_fill_1 FILLER_20_128 ();
 sg13g2_fill_1 FILLER_20_142 ();
 sg13g2_fill_1 FILLER_20_150 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_4 FILLER_20_179 ();
 sg13g2_fill_1 FILLER_20_183 ();
 sg13g2_decap_4 FILLER_20_197 ();
 sg13g2_fill_1 FILLER_20_201 ();
 sg13g2_decap_4 FILLER_20_215 ();
 sg13g2_decap_4 FILLER_20_233 ();
 sg13g2_fill_1 FILLER_20_237 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_fill_2 FILLER_20_284 ();
 sg13g2_fill_1 FILLER_20_286 ();
 sg13g2_fill_2 FILLER_20_300 ();
 sg13g2_fill_1 FILLER_20_307 ();
 sg13g2_fill_1 FILLER_20_314 ();
 sg13g2_fill_1 FILLER_20_337 ();
 sg13g2_decap_8 FILLER_20_364 ();
 sg13g2_decap_8 FILLER_20_371 ();
 sg13g2_decap_8 FILLER_20_378 ();
 sg13g2_decap_8 FILLER_20_385 ();
 sg13g2_decap_8 FILLER_20_392 ();
 sg13g2_decap_8 FILLER_20_399 ();
 sg13g2_fill_2 FILLER_20_406 ();
 sg13g2_fill_1 FILLER_20_408 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_fill_2 FILLER_21_14 ();
 sg13g2_fill_2 FILLER_21_29 ();
 sg13g2_fill_2 FILLER_21_36 ();
 sg13g2_fill_1 FILLER_21_38 ();
 sg13g2_fill_2 FILLER_21_52 ();
 sg13g2_fill_1 FILLER_21_54 ();
 sg13g2_decap_8 FILLER_21_69 ();
 sg13g2_decap_8 FILLER_21_76 ();
 sg13g2_decap_8 FILLER_21_83 ();
 sg13g2_fill_1 FILLER_21_90 ();
 sg13g2_decap_8 FILLER_21_99 ();
 sg13g2_decap_8 FILLER_21_106 ();
 sg13g2_fill_1 FILLER_21_113 ();
 sg13g2_decap_8 FILLER_21_127 ();
 sg13g2_decap_4 FILLER_21_134 ();
 sg13g2_fill_2 FILLER_21_156 ();
 sg13g2_fill_1 FILLER_21_158 ();
 sg13g2_decap_4 FILLER_21_173 ();
 sg13g2_fill_1 FILLER_21_184 ();
 sg13g2_decap_4 FILLER_21_198 ();
 sg13g2_fill_1 FILLER_21_209 ();
 sg13g2_decap_8 FILLER_21_237 ();
 sg13g2_decap_4 FILLER_21_244 ();
 sg13g2_fill_2 FILLER_21_248 ();
 sg13g2_fill_2 FILLER_21_255 ();
 sg13g2_fill_2 FILLER_21_261 ();
 sg13g2_fill_1 FILLER_21_263 ();
 sg13g2_decap_8 FILLER_21_270 ();
 sg13g2_decap_8 FILLER_21_277 ();
 sg13g2_fill_2 FILLER_21_284 ();
 sg13g2_fill_1 FILLER_21_286 ();
 sg13g2_fill_2 FILLER_21_335 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_fill_2 FILLER_21_406 ();
 sg13g2_fill_1 FILLER_21_408 ();
 sg13g2_decap_8 FILLER_22_0 ();
 sg13g2_decap_8 FILLER_22_7 ();
 sg13g2_decap_8 FILLER_22_14 ();
 sg13g2_decap_8 FILLER_22_21 ();
 sg13g2_fill_2 FILLER_22_28 ();
 sg13g2_fill_1 FILLER_22_30 ();
 sg13g2_fill_1 FILLER_22_46 ();
 sg13g2_fill_1 FILLER_22_66 ();
 sg13g2_fill_1 FILLER_22_77 ();
 sg13g2_decap_4 FILLER_22_103 ();
 sg13g2_fill_2 FILLER_22_145 ();
 sg13g2_decap_8 FILLER_22_157 ();
 sg13g2_decap_8 FILLER_22_164 ();
 sg13g2_fill_2 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_246 ();
 sg13g2_decap_8 FILLER_22_253 ();
 sg13g2_decap_4 FILLER_22_260 ();
 sg13g2_decap_8 FILLER_22_272 ();
 sg13g2_decap_4 FILLER_22_279 ();
 sg13g2_fill_1 FILLER_22_283 ();
 sg13g2_fill_2 FILLER_22_314 ();
 sg13g2_fill_2 FILLER_22_327 ();
 sg13g2_fill_1 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_4 FILLER_22_403 ();
 sg13g2_fill_2 FILLER_22_407 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_fill_1 FILLER_23_45 ();
 sg13g2_fill_2 FILLER_23_135 ();
 sg13g2_fill_1 FILLER_23_137 ();
 sg13g2_decap_8 FILLER_23_162 ();
 sg13g2_decap_8 FILLER_23_169 ();
 sg13g2_fill_1 FILLER_23_176 ();
 sg13g2_fill_2 FILLER_23_181 ();
 sg13g2_decap_8 FILLER_23_206 ();
 sg13g2_fill_2 FILLER_23_225 ();
 sg13g2_fill_1 FILLER_23_227 ();
 sg13g2_fill_2 FILLER_23_233 ();
 sg13g2_fill_1 FILLER_23_235 ();
 sg13g2_decap_8 FILLER_23_264 ();
 sg13g2_decap_4 FILLER_23_271 ();
 sg13g2_decap_8 FILLER_23_281 ();
 sg13g2_decap_8 FILLER_23_288 ();
 sg13g2_decap_8 FILLER_23_295 ();
 sg13g2_fill_2 FILLER_23_302 ();
 sg13g2_fill_1 FILLER_23_304 ();
 sg13g2_fill_2 FILLER_23_349 ();
 sg13g2_decap_4 FILLER_23_356 ();
 sg13g2_fill_1 FILLER_23_360 ();
 sg13g2_decap_8 FILLER_23_366 ();
 sg13g2_decap_8 FILLER_23_373 ();
 sg13g2_decap_8 FILLER_23_380 ();
 sg13g2_decap_8 FILLER_23_387 ();
 sg13g2_decap_8 FILLER_23_394 ();
 sg13g2_decap_8 FILLER_23_401 ();
 sg13g2_fill_1 FILLER_23_408 ();
 sg13g2_decap_8 FILLER_24_0 ();
 sg13g2_decap_8 FILLER_24_7 ();
 sg13g2_decap_8 FILLER_24_14 ();
 sg13g2_fill_2 FILLER_24_21 ();
 sg13g2_fill_2 FILLER_24_31 ();
 sg13g2_fill_1 FILLER_24_33 ();
 sg13g2_fill_1 FILLER_24_38 ();
 sg13g2_decap_8 FILLER_24_52 ();
 sg13g2_fill_1 FILLER_24_59 ();
 sg13g2_decap_8 FILLER_24_82 ();
 sg13g2_decap_8 FILLER_24_101 ();
 sg13g2_decap_4 FILLER_24_108 ();
 sg13g2_fill_2 FILLER_24_112 ();
 sg13g2_fill_1 FILLER_24_131 ();
 sg13g2_fill_1 FILLER_24_148 ();
 sg13g2_fill_1 FILLER_24_154 ();
 sg13g2_fill_2 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_171 ();
 sg13g2_decap_8 FILLER_24_178 ();
 sg13g2_decap_4 FILLER_24_185 ();
 sg13g2_decap_4 FILLER_24_197 ();
 sg13g2_fill_2 FILLER_24_201 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_fill_1 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_280 ();
 sg13g2_fill_2 FILLER_24_287 ();
 sg13g2_fill_2 FILLER_24_294 ();
 sg13g2_decap_8 FILLER_24_307 ();
 sg13g2_decap_8 FILLER_24_314 ();
 sg13g2_fill_1 FILLER_24_321 ();
 sg13g2_decap_4 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_348 ();
 sg13g2_fill_2 FILLER_24_355 ();
 sg13g2_fill_1 FILLER_24_357 ();
 sg13g2_fill_1 FILLER_24_362 ();
 sg13g2_decap_8 FILLER_24_367 ();
 sg13g2_decap_8 FILLER_24_374 ();
 sg13g2_decap_8 FILLER_24_381 ();
 sg13g2_decap_8 FILLER_24_388 ();
 sg13g2_decap_8 FILLER_24_395 ();
 sg13g2_decap_8 FILLER_24_402 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_fill_1 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_58 ();
 sg13g2_decap_8 FILLER_25_65 ();
 sg13g2_decap_8 FILLER_25_72 ();
 sg13g2_decap_8 FILLER_25_79 ();
 sg13g2_decap_8 FILLER_25_100 ();
 sg13g2_decap_8 FILLER_25_107 ();
 sg13g2_decap_4 FILLER_25_114 ();
 sg13g2_fill_2 FILLER_25_118 ();
 sg13g2_fill_2 FILLER_25_177 ();
 sg13g2_fill_1 FILLER_25_179 ();
 sg13g2_fill_2 FILLER_25_189 ();
 sg13g2_fill_1 FILLER_25_191 ();
 sg13g2_fill_2 FILLER_25_255 ();
 sg13g2_fill_1 FILLER_25_270 ();
 sg13g2_fill_2 FILLER_25_276 ();
 sg13g2_decap_4 FILLER_25_284 ();
 sg13g2_fill_1 FILLER_25_297 ();
 sg13g2_fill_2 FILLER_25_311 ();
 sg13g2_fill_2 FILLER_25_325 ();
 sg13g2_fill_1 FILLER_25_327 ();
 sg13g2_decap_8 FILLER_25_333 ();
 sg13g2_decap_8 FILLER_25_340 ();
 sg13g2_fill_2 FILLER_25_368 ();
 sg13g2_fill_1 FILLER_25_370 ();
 sg13g2_decap_8 FILLER_25_379 ();
 sg13g2_decap_8 FILLER_25_386 ();
 sg13g2_decap_8 FILLER_25_393 ();
 sg13g2_decap_8 FILLER_25_400 ();
 sg13g2_fill_2 FILLER_25_407 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_fill_1 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_13 ();
 sg13g2_decap_8 FILLER_26_30 ();
 sg13g2_fill_2 FILLER_26_37 ();
 sg13g2_decap_8 FILLER_26_52 ();
 sg13g2_decap_8 FILLER_26_59 ();
 sg13g2_decap_8 FILLER_26_66 ();
 sg13g2_fill_2 FILLER_26_73 ();
 sg13g2_fill_1 FILLER_26_75 ();
 sg13g2_fill_1 FILLER_26_103 ();
 sg13g2_decap_4 FILLER_26_108 ();
 sg13g2_fill_2 FILLER_26_112 ();
 sg13g2_fill_2 FILLER_26_121 ();
 sg13g2_fill_2 FILLER_26_141 ();
 sg13g2_fill_1 FILLER_26_143 ();
 sg13g2_fill_2 FILLER_26_152 ();
 sg13g2_fill_1 FILLER_26_154 ();
 sg13g2_fill_1 FILLER_26_163 ();
 sg13g2_fill_2 FILLER_26_172 ();
 sg13g2_fill_2 FILLER_26_182 ();
 sg13g2_fill_1 FILLER_26_184 ();
 sg13g2_fill_2 FILLER_26_197 ();
 sg13g2_fill_2 FILLER_26_237 ();
 sg13g2_decap_4 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_270 ();
 sg13g2_fill_1 FILLER_26_291 ();
 sg13g2_decap_4 FILLER_26_297 ();
 sg13g2_decap_8 FILLER_26_321 ();
 sg13g2_decap_4 FILLER_26_350 ();
 sg13g2_fill_2 FILLER_26_359 ();
 sg13g2_fill_1 FILLER_26_361 ();
 sg13g2_fill_2 FILLER_26_367 ();
 sg13g2_decap_8 FILLER_26_374 ();
 sg13g2_decap_8 FILLER_26_381 ();
 sg13g2_decap_8 FILLER_26_388 ();
 sg13g2_decap_8 FILLER_26_395 ();
 sg13g2_decap_8 FILLER_26_402 ();
 sg13g2_fill_2 FILLER_27_0 ();
 sg13g2_fill_1 FILLER_27_2 ();
 sg13g2_decap_4 FILLER_27_24 ();
 sg13g2_fill_2 FILLER_27_28 ();
 sg13g2_fill_2 FILLER_27_35 ();
 sg13g2_fill_2 FILLER_27_50 ();
 sg13g2_fill_1 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_152 ();
 sg13g2_fill_2 FILLER_27_159 ();
 sg13g2_fill_1 FILLER_27_161 ();
 sg13g2_fill_1 FILLER_27_182 ();
 sg13g2_fill_1 FILLER_27_201 ();
 sg13g2_fill_2 FILLER_27_207 ();
 sg13g2_fill_1 FILLER_27_217 ();
 sg13g2_decap_8 FILLER_27_227 ();
 sg13g2_decap_4 FILLER_27_234 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_4 FILLER_27_249 ();
 sg13g2_fill_2 FILLER_27_253 ();
 sg13g2_decap_8 FILLER_27_260 ();
 sg13g2_decap_4 FILLER_27_267 ();
 sg13g2_fill_2 FILLER_27_271 ();
 sg13g2_decap_4 FILLER_27_280 ();
 sg13g2_fill_2 FILLER_27_284 ();
 sg13g2_fill_2 FILLER_27_298 ();
 sg13g2_fill_1 FILLER_27_300 ();
 sg13g2_decap_4 FILLER_27_307 ();
 sg13g2_fill_1 FILLER_27_311 ();
 sg13g2_decap_4 FILLER_27_342 ();
 sg13g2_fill_1 FILLER_27_346 ();
 sg13g2_decap_8 FILLER_27_387 ();
 sg13g2_decap_8 FILLER_27_394 ();
 sg13g2_decap_8 FILLER_27_401 ();
 sg13g2_fill_1 FILLER_27_408 ();
 sg13g2_decap_4 FILLER_28_0 ();
 sg13g2_fill_2 FILLER_28_60 ();
 sg13g2_fill_1 FILLER_28_62 ();
 sg13g2_decap_4 FILLER_28_133 ();
 sg13g2_decap_4 FILLER_28_155 ();
 sg13g2_decap_4 FILLER_28_165 ();
 sg13g2_fill_2 FILLER_28_174 ();
 sg13g2_fill_1 FILLER_28_176 ();
 sg13g2_fill_2 FILLER_28_187 ();
 sg13g2_fill_1 FILLER_28_189 ();
 sg13g2_decap_4 FILLER_28_224 ();
 sg13g2_fill_2 FILLER_28_228 ();
 sg13g2_fill_2 FILLER_28_235 ();
 sg13g2_fill_1 FILLER_28_237 ();
 sg13g2_fill_2 FILLER_28_243 ();
 sg13g2_fill_1 FILLER_28_268 ();
 sg13g2_decap_4 FILLER_28_285 ();
 sg13g2_fill_1 FILLER_28_289 ();
 sg13g2_fill_2 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_321 ();
 sg13g2_decap_4 FILLER_28_328 ();
 sg13g2_decap_8 FILLER_28_342 ();
 sg13g2_decap_8 FILLER_28_349 ();
 sg13g2_fill_1 FILLER_28_356 ();
 sg13g2_decap_8 FILLER_28_363 ();
 sg13g2_decap_4 FILLER_28_370 ();
 sg13g2_fill_1 FILLER_28_374 ();
 sg13g2_decap_8 FILLER_28_381 ();
 sg13g2_decap_8 FILLER_28_388 ();
 sg13g2_decap_8 FILLER_28_395 ();
 sg13g2_decap_8 FILLER_28_402 ();
 sg13g2_fill_2 FILLER_29_0 ();
 sg13g2_fill_1 FILLER_29_2 ();
 sg13g2_fill_2 FILLER_29_36 ();
 sg13g2_decap_8 FILLER_29_51 ();
 sg13g2_fill_1 FILLER_29_58 ();
 sg13g2_decap_8 FILLER_29_73 ();
 sg13g2_decap_4 FILLER_29_80 ();
 sg13g2_fill_1 FILLER_29_84 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_fill_1 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_143 ();
 sg13g2_decap_8 FILLER_29_150 ();
 sg13g2_decap_4 FILLER_29_174 ();
 sg13g2_decap_4 FILLER_29_183 ();
 sg13g2_fill_2 FILLER_29_187 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_fill_1 FILLER_29_200 ();
 sg13g2_decap_4 FILLER_29_209 ();
 sg13g2_fill_2 FILLER_29_213 ();
 sg13g2_fill_1 FILLER_29_253 ();
 sg13g2_fill_1 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_282 ();
 sg13g2_decap_4 FILLER_29_289 ();
 sg13g2_fill_2 FILLER_29_293 ();
 sg13g2_decap_8 FILLER_29_310 ();
 sg13g2_decap_8 FILLER_29_317 ();
 sg13g2_fill_1 FILLER_29_328 ();
 sg13g2_fill_2 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_fill_2 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_369 ();
 sg13g2_decap_8 FILLER_29_376 ();
 sg13g2_decap_8 FILLER_29_383 ();
 sg13g2_decap_8 FILLER_29_390 ();
 sg13g2_decap_8 FILLER_29_397 ();
 sg13g2_decap_4 FILLER_29_404 ();
 sg13g2_fill_1 FILLER_29_408 ();
 sg13g2_decap_4 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_38 ();
 sg13g2_decap_8 FILLER_30_45 ();
 sg13g2_fill_2 FILLER_30_52 ();
 sg13g2_decap_4 FILLER_30_68 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_fill_2 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_fill_2 FILLER_30_112 ();
 sg13g2_fill_1 FILLER_30_114 ();
 sg13g2_decap_4 FILLER_30_120 ();
 sg13g2_fill_2 FILLER_30_124 ();
 sg13g2_decap_8 FILLER_30_134 ();
 sg13g2_decap_8 FILLER_30_141 ();
 sg13g2_decap_8 FILLER_30_169 ();
 sg13g2_decap_4 FILLER_30_176 ();
 sg13g2_fill_2 FILLER_30_180 ();
 sg13g2_fill_1 FILLER_30_188 ();
 sg13g2_decap_4 FILLER_30_202 ();
 sg13g2_fill_1 FILLER_30_206 ();
 sg13g2_fill_2 FILLER_30_260 ();
 sg13g2_fill_1 FILLER_30_262 ();
 sg13g2_decap_8 FILLER_30_268 ();
 sg13g2_decap_8 FILLER_30_275 ();
 sg13g2_decap_8 FILLER_30_282 ();
 sg13g2_fill_1 FILLER_30_289 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_fill_2 FILLER_30_308 ();
 sg13g2_fill_1 FILLER_30_310 ();
 sg13g2_fill_2 FILLER_30_320 ();
 sg13g2_fill_1 FILLER_30_322 ();
 sg13g2_fill_2 FILLER_30_352 ();
 sg13g2_fill_1 FILLER_30_354 ();
 sg13g2_fill_2 FILLER_30_360 ();
 sg13g2_fill_1 FILLER_30_362 ();
 sg13g2_fill_2 FILLER_30_372 ();
 sg13g2_decap_8 FILLER_30_379 ();
 sg13g2_decap_8 FILLER_30_386 ();
 sg13g2_decap_8 FILLER_30_393 ();
 sg13g2_decap_8 FILLER_30_400 ();
 sg13g2_fill_2 FILLER_30_407 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_fill_1 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_25 ();
 sg13g2_decap_8 FILLER_31_32 ();
 sg13g2_decap_8 FILLER_31_39 ();
 sg13g2_decap_8 FILLER_31_46 ();
 sg13g2_fill_2 FILLER_31_53 ();
 sg13g2_fill_1 FILLER_31_55 ();
 sg13g2_fill_2 FILLER_31_62 ();
 sg13g2_fill_2 FILLER_31_72 ();
 sg13g2_decap_8 FILLER_31_80 ();
 sg13g2_decap_8 FILLER_31_95 ();
 sg13g2_decap_8 FILLER_31_102 ();
 sg13g2_fill_2 FILLER_31_177 ();
 sg13g2_fill_1 FILLER_31_179 ();
 sg13g2_fill_2 FILLER_31_202 ();
 sg13g2_fill_1 FILLER_31_204 ();
 sg13g2_fill_2 FILLER_31_257 ();
 sg13g2_fill_1 FILLER_31_259 ();
 sg13g2_decap_4 FILLER_31_291 ();
 sg13g2_fill_2 FILLER_31_295 ();
 sg13g2_fill_2 FILLER_31_324 ();
 sg13g2_decap_8 FILLER_31_347 ();
 sg13g2_decap_8 FILLER_31_354 ();
 sg13g2_decap_8 FILLER_31_361 ();
 sg13g2_decap_4 FILLER_31_368 ();
 sg13g2_fill_1 FILLER_31_372 ();
 sg13g2_decap_8 FILLER_31_387 ();
 sg13g2_decap_8 FILLER_31_394 ();
 sg13g2_decap_8 FILLER_31_401 ();
 sg13g2_fill_1 FILLER_31_408 ();
 sg13g2_decap_4 FILLER_32_0 ();
 sg13g2_fill_1 FILLER_32_4 ();
 sg13g2_fill_1 FILLER_32_30 ();
 sg13g2_fill_1 FILLER_32_43 ();
 sg13g2_decap_4 FILLER_32_49 ();
 sg13g2_fill_1 FILLER_32_69 ();
 sg13g2_decap_4 FILLER_32_94 ();
 sg13g2_fill_2 FILLER_32_98 ();
 sg13g2_fill_1 FILLER_32_138 ();
 sg13g2_fill_2 FILLER_32_147 ();
 sg13g2_decap_8 FILLER_32_169 ();
 sg13g2_fill_2 FILLER_32_176 ();
 sg13g2_fill_1 FILLER_32_178 ();
 sg13g2_fill_1 FILLER_32_211 ();
 sg13g2_decap_4 FILLER_32_248 ();
 sg13g2_fill_2 FILLER_32_252 ();
 sg13g2_decap_4 FILLER_32_258 ();
 sg13g2_fill_2 FILLER_32_268 ();
 sg13g2_fill_1 FILLER_32_270 ();
 sg13g2_decap_4 FILLER_32_284 ();
 sg13g2_fill_1 FILLER_32_306 ();
 sg13g2_fill_2 FILLER_32_316 ();
 sg13g2_fill_1 FILLER_32_318 ();
 sg13g2_fill_1 FILLER_32_324 ();
 sg13g2_decap_4 FILLER_32_333 ();
 sg13g2_fill_1 FILLER_32_337 ();
 sg13g2_fill_1 FILLER_32_342 ();
 sg13g2_decap_4 FILLER_32_349 ();
 sg13g2_fill_1 FILLER_32_353 ();
 sg13g2_decap_4 FILLER_32_364 ();
 sg13g2_decap_8 FILLER_32_373 ();
 sg13g2_decap_8 FILLER_32_380 ();
 sg13g2_decap_8 FILLER_32_387 ();
 sg13g2_decap_8 FILLER_32_394 ();
 sg13g2_decap_8 FILLER_32_401 ();
 sg13g2_fill_1 FILLER_32_408 ();
 sg13g2_fill_2 FILLER_33_0 ();
 sg13g2_fill_1 FILLER_33_25 ();
 sg13g2_fill_1 FILLER_33_60 ();
 sg13g2_fill_2 FILLER_33_95 ();
 sg13g2_fill_1 FILLER_33_97 ();
 sg13g2_fill_2 FILLER_33_110 ();
 sg13g2_fill_1 FILLER_33_112 ();
 sg13g2_fill_2 FILLER_33_132 ();
 sg13g2_decap_4 FILLER_33_147 ();
 sg13g2_fill_1 FILLER_33_151 ();
 sg13g2_decap_4 FILLER_33_157 ();
 sg13g2_fill_2 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_4 FILLER_33_182 ();
 sg13g2_fill_2 FILLER_33_186 ();
 sg13g2_fill_1 FILLER_33_196 ();
 sg13g2_fill_2 FILLER_33_205 ();
 sg13g2_decap_8 FILLER_33_213 ();
 sg13g2_decap_8 FILLER_33_220 ();
 sg13g2_decap_8 FILLER_33_227 ();
 sg13g2_fill_2 FILLER_33_234 ();
 sg13g2_decap_8 FILLER_33_244 ();
 sg13g2_decap_4 FILLER_33_251 ();
 sg13g2_fill_2 FILLER_33_255 ();
 sg13g2_decap_4 FILLER_33_261 ();
 sg13g2_fill_1 FILLER_33_265 ();
 sg13g2_fill_2 FILLER_33_285 ();
 sg13g2_decap_8 FILLER_33_302 ();
 sg13g2_decap_8 FILLER_33_313 ();
 sg13g2_decap_4 FILLER_33_320 ();
 sg13g2_decap_4 FILLER_33_329 ();
 sg13g2_fill_1 FILLER_33_333 ();
 sg13g2_decap_8 FILLER_33_339 ();
 sg13g2_decap_4 FILLER_33_346 ();
 sg13g2_decap_4 FILLER_33_355 ();
 sg13g2_fill_2 FILLER_33_359 ();
 sg13g2_decap_8 FILLER_33_374 ();
 sg13g2_decap_8 FILLER_33_381 ();
 sg13g2_decap_8 FILLER_33_388 ();
 sg13g2_decap_8 FILLER_33_395 ();
 sg13g2_decap_8 FILLER_33_402 ();
 sg13g2_fill_2 FILLER_34_0 ();
 sg13g2_fill_1 FILLER_34_2 ();
 sg13g2_fill_2 FILLER_34_33 ();
 sg13g2_decap_4 FILLER_34_45 ();
 sg13g2_fill_1 FILLER_34_49 ();
 sg13g2_decap_8 FILLER_34_63 ();
 sg13g2_fill_2 FILLER_34_70 ();
 sg13g2_fill_1 FILLER_34_72 ();
 sg13g2_fill_2 FILLER_34_78 ();
 sg13g2_fill_1 FILLER_34_80 ();
 sg13g2_decap_4 FILLER_34_105 ();
 sg13g2_decap_4 FILLER_34_124 ();
 sg13g2_fill_2 FILLER_34_128 ();
 sg13g2_fill_2 FILLER_34_134 ();
 sg13g2_fill_1 FILLER_34_136 ();
 sg13g2_decap_8 FILLER_34_141 ();
 sg13g2_fill_2 FILLER_34_148 ();
 sg13g2_decap_8 FILLER_34_176 ();
 sg13g2_decap_8 FILLER_34_183 ();
 sg13g2_decap_4 FILLER_34_190 ();
 sg13g2_decap_8 FILLER_34_199 ();
 sg13g2_decap_4 FILLER_34_206 ();
 sg13g2_fill_1 FILLER_34_210 ();
 sg13g2_fill_2 FILLER_34_225 ();
 sg13g2_decap_4 FILLER_34_236 ();
 sg13g2_fill_1 FILLER_34_240 ();
 sg13g2_fill_1 FILLER_34_275 ();
 sg13g2_decap_8 FILLER_34_296 ();
 sg13g2_decap_8 FILLER_34_303 ();
 sg13g2_decap_4 FILLER_34_310 ();
 sg13g2_decap_8 FILLER_34_350 ();
 sg13g2_decap_8 FILLER_34_357 ();
 sg13g2_decap_8 FILLER_34_364 ();
 sg13g2_decap_8 FILLER_34_371 ();
 sg13g2_decap_4 FILLER_34_378 ();
 sg13g2_fill_2 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_395 ();
 sg13g2_decap_8 FILLER_34_402 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_fill_2 FILLER_35_14 ();
 sg13g2_fill_1 FILLER_35_16 ();
 sg13g2_fill_2 FILLER_35_22 ();
 sg13g2_fill_1 FILLER_35_24 ();
 sg13g2_decap_8 FILLER_35_31 ();
 sg13g2_decap_8 FILLER_35_38 ();
 sg13g2_decap_8 FILLER_35_45 ();
 sg13g2_decap_8 FILLER_35_52 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_fill_2 FILLER_35_98 ();
 sg13g2_fill_1 FILLER_35_100 ();
 sg13g2_fill_2 FILLER_35_107 ();
 sg13g2_fill_1 FILLER_35_109 ();
 sg13g2_decap_4 FILLER_35_148 ();
 sg13g2_fill_2 FILLER_35_152 ();
 sg13g2_fill_1 FILLER_35_180 ();
 sg13g2_decap_8 FILLER_35_187 ();
 sg13g2_decap_8 FILLER_35_194 ();
 sg13g2_decap_4 FILLER_35_201 ();
 sg13g2_fill_1 FILLER_35_205 ();
 sg13g2_fill_2 FILLER_35_234 ();
 sg13g2_fill_1 FILLER_35_236 ();
 sg13g2_fill_2 FILLER_35_250 ();
 sg13g2_fill_1 FILLER_35_252 ();
 sg13g2_fill_1 FILLER_35_284 ();
 sg13g2_fill_1 FILLER_35_304 ();
 sg13g2_decap_4 FILLER_35_313 ();
 sg13g2_fill_2 FILLER_35_317 ();
 sg13g2_decap_8 FILLER_35_335 ();
 sg13g2_fill_2 FILLER_35_342 ();
 sg13g2_fill_1 FILLER_35_344 ();
 sg13g2_decap_8 FILLER_35_358 ();
 sg13g2_decap_8 FILLER_35_365 ();
 sg13g2_decap_8 FILLER_35_376 ();
 sg13g2_fill_2 FILLER_35_383 ();
 sg13g2_fill_1 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_396 ();
 sg13g2_decap_4 FILLER_35_403 ();
 sg13g2_fill_2 FILLER_35_407 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_fill_1 FILLER_36_21 ();
 sg13g2_decap_4 FILLER_36_26 ();
 sg13g2_fill_2 FILLER_36_30 ();
 sg13g2_fill_2 FILLER_36_37 ();
 sg13g2_fill_1 FILLER_36_39 ();
 sg13g2_fill_1 FILLER_36_45 ();
 sg13g2_decap_8 FILLER_36_76 ();
 sg13g2_fill_1 FILLER_36_93 ();
 sg13g2_fill_1 FILLER_36_107 ();
 sg13g2_fill_2 FILLER_36_127 ();
 sg13g2_decap_8 FILLER_36_153 ();
 sg13g2_fill_2 FILLER_36_160 ();
 sg13g2_fill_1 FILLER_36_186 ();
 sg13g2_fill_2 FILLER_36_208 ();
 sg13g2_fill_2 FILLER_36_223 ();
 sg13g2_fill_1 FILLER_36_225 ();
 sg13g2_fill_1 FILLER_36_235 ();
 sg13g2_fill_1 FILLER_36_253 ();
 sg13g2_fill_2 FILLER_36_259 ();
 sg13g2_fill_1 FILLER_36_303 ();
 sg13g2_decap_8 FILLER_36_320 ();
 sg13g2_decap_4 FILLER_36_327 ();
 sg13g2_fill_1 FILLER_36_331 ();
 sg13g2_decap_4 FILLER_36_338 ();
 sg13g2_fill_2 FILLER_36_342 ();
 sg13g2_decap_4 FILLER_36_348 ();
 sg13g2_fill_2 FILLER_36_352 ();
 sg13g2_fill_2 FILLER_36_364 ();
 sg13g2_fill_1 FILLER_36_366 ();
 sg13g2_fill_2 FILLER_36_377 ();
 sg13g2_decap_4 FILLER_36_403 ();
 sg13g2_fill_2 FILLER_36_407 ();
 sg13g2_decap_8 FILLER_37_0 ();
 sg13g2_fill_2 FILLER_37_20 ();
 sg13g2_fill_1 FILLER_37_22 ();
 sg13g2_fill_1 FILLER_37_55 ();
 sg13g2_fill_2 FILLER_37_70 ();
 sg13g2_fill_1 FILLER_37_72 ();
 sg13g2_fill_2 FILLER_37_81 ();
 sg13g2_fill_2 FILLER_37_101 ();
 sg13g2_fill_1 FILLER_37_103 ();
 sg13g2_fill_1 FILLER_37_127 ();
 sg13g2_decap_4 FILLER_37_172 ();
 sg13g2_decap_4 FILLER_37_180 ();
 sg13g2_fill_2 FILLER_37_184 ();
 sg13g2_fill_1 FILLER_37_199 ();
 sg13g2_fill_1 FILLER_37_213 ();
 sg13g2_fill_1 FILLER_37_218 ();
 sg13g2_fill_2 FILLER_37_251 ();
 sg13g2_fill_1 FILLER_37_253 ();
 sg13g2_decap_4 FILLER_37_264 ();
 sg13g2_fill_2 FILLER_37_281 ();
 sg13g2_fill_1 FILLER_37_289 ();
 sg13g2_decap_4 FILLER_37_308 ();
 sg13g2_decap_4 FILLER_37_318 ();
 sg13g2_fill_2 FILLER_37_322 ();
 sg13g2_decap_4 FILLER_37_330 ();
 sg13g2_fill_1 FILLER_37_334 ();
 sg13g2_fill_1 FILLER_37_346 ();
 sg13g2_fill_1 FILLER_37_356 ();
 sg13g2_decap_8 FILLER_37_376 ();
 sg13g2_decap_4 FILLER_37_383 ();
 sg13g2_fill_2 FILLER_37_393 ();
 sg13g2_fill_1 FILLER_37_395 ();
 sg13g2_fill_2 FILLER_37_407 ();
 sg13g2_fill_2 FILLER_38_0 ();
 sg13g2_fill_1 FILLER_38_2 ();
 sg13g2_fill_1 FILLER_38_29 ();
 sg13g2_fill_2 FILLER_38_62 ();
 sg13g2_fill_1 FILLER_38_88 ();
 sg13g2_fill_1 FILLER_38_119 ();
 sg13g2_fill_1 FILLER_38_143 ();
 sg13g2_fill_1 FILLER_38_154 ();
 sg13g2_fill_2 FILLER_38_173 ();
 sg13g2_fill_1 FILLER_38_175 ();
 sg13g2_fill_1 FILLER_38_228 ();
 sg13g2_fill_2 FILLER_38_243 ();
 sg13g2_fill_1 FILLER_38_249 ();
 sg13g2_decap_8 FILLER_38_260 ();
 sg13g2_fill_2 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_306 ();
 sg13g2_fill_1 FILLER_38_313 ();
 sg13g2_decap_8 FILLER_38_338 ();
 sg13g2_decap_8 FILLER_38_345 ();
 sg13g2_decap_4 FILLER_38_352 ();
 sg13g2_fill_1 FILLER_38_365 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_fill_2 FILLER_38_406 ();
 sg13g2_fill_1 FILLER_38_408 ();
 sg13g2_fill_2 FILLER_39_0 ();
 sg13g2_fill_1 FILLER_39_2 ();
 sg13g2_decap_4 FILLER_39_21 ();
 sg13g2_fill_2 FILLER_39_43 ();
 sg13g2_fill_1 FILLER_39_45 ();
 sg13g2_fill_1 FILLER_39_59 ();
 sg13g2_fill_1 FILLER_39_92 ();
 sg13g2_decap_4 FILLER_39_112 ();
 sg13g2_fill_1 FILLER_39_116 ();
 sg13g2_fill_2 FILLER_39_127 ();
 sg13g2_fill_1 FILLER_39_129 ();
 sg13g2_fill_2 FILLER_39_146 ();
 sg13g2_fill_2 FILLER_39_154 ();
 sg13g2_fill_2 FILLER_39_182 ();
 sg13g2_decap_8 FILLER_39_189 ();
 sg13g2_decap_4 FILLER_39_196 ();
 sg13g2_fill_1 FILLER_39_200 ();
 sg13g2_decap_4 FILLER_39_207 ();
 sg13g2_fill_2 FILLER_39_260 ();
 sg13g2_fill_2 FILLER_39_270 ();
 sg13g2_fill_2 FILLER_39_282 ();
 sg13g2_fill_2 FILLER_39_290 ();
 sg13g2_fill_1 FILLER_39_292 ();
 sg13g2_fill_2 FILLER_39_299 ();
 sg13g2_fill_1 FILLER_39_301 ();
 sg13g2_fill_1 FILLER_39_314 ();
 sg13g2_decap_4 FILLER_39_320 ();
 sg13g2_fill_2 FILLER_39_324 ();
 sg13g2_decap_8 FILLER_39_341 ();
 sg13g2_decap_8 FILLER_39_348 ();
 sg13g2_decap_8 FILLER_39_355 ();
 sg13g2_fill_1 FILLER_39_362 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_decap_4 FILLER_39_389 ();
 sg13g2_fill_2 FILLER_39_393 ();
 sg13g2_decap_8 FILLER_39_400 ();
 sg13g2_fill_2 FILLER_39_407 ();
 sg13g2_fill_1 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_19 ();
 sg13g2_decap_8 FILLER_40_26 ();
 sg13g2_decap_8 FILLER_40_33 ();
 sg13g2_fill_1 FILLER_40_40 ();
 sg13g2_decap_8 FILLER_40_46 ();
 sg13g2_decap_8 FILLER_40_53 ();
 sg13g2_decap_4 FILLER_40_60 ();
 sg13g2_fill_1 FILLER_40_64 ();
 sg13g2_decap_8 FILLER_40_76 ();
 sg13g2_decap_8 FILLER_40_83 ();
 sg13g2_decap_4 FILLER_40_90 ();
 sg13g2_fill_2 FILLER_40_94 ();
 sg13g2_decap_8 FILLER_40_101 ();
 sg13g2_decap_4 FILLER_40_108 ();
 sg13g2_fill_2 FILLER_40_125 ();
 sg13g2_fill_2 FILLER_40_145 ();
 sg13g2_fill_1 FILLER_40_147 ();
 sg13g2_decap_4 FILLER_40_152 ();
 sg13g2_fill_1 FILLER_40_156 ();
 sg13g2_decap_8 FILLER_40_162 ();
 sg13g2_fill_1 FILLER_40_169 ();
 sg13g2_fill_1 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_181 ();
 sg13g2_decap_4 FILLER_40_188 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_4 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_226 ();
 sg13g2_fill_2 FILLER_40_233 ();
 sg13g2_fill_1 FILLER_40_235 ();
 sg13g2_fill_2 FILLER_40_246 ();
 sg13g2_fill_2 FILLER_40_267 ();
 sg13g2_fill_2 FILLER_40_279 ();
 sg13g2_fill_1 FILLER_40_294 ();
 sg13g2_fill_2 FILLER_40_314 ();
 sg13g2_fill_1 FILLER_40_316 ();
 sg13g2_fill_2 FILLER_40_323 ();
 sg13g2_fill_1 FILLER_40_325 ();
 sg13g2_fill_1 FILLER_40_342 ();
 sg13g2_decap_8 FILLER_40_354 ();
 sg13g2_fill_2 FILLER_40_361 ();
 sg13g2_fill_1 FILLER_40_363 ();
 sg13g2_decap_4 FILLER_40_372 ();
 sg13g2_fill_2 FILLER_40_376 ();
 sg13g2_decap_8 FILLER_40_395 ();
 sg13g2_decap_8 FILLER_40_402 ();
 sg13g2_decap_4 FILLER_41_0 ();
 sg13g2_fill_1 FILLER_41_25 ();
 sg13g2_decap_8 FILLER_41_68 ();
 sg13g2_fill_2 FILLER_41_75 ();
 sg13g2_fill_1 FILLER_41_77 ();
 sg13g2_fill_2 FILLER_41_93 ();
 sg13g2_fill_1 FILLER_41_95 ();
 sg13g2_decap_4 FILLER_41_101 ();
 sg13g2_fill_2 FILLER_41_105 ();
 sg13g2_fill_1 FILLER_41_133 ();
 sg13g2_fill_1 FILLER_41_140 ();
 sg13g2_fill_2 FILLER_41_153 ();
 sg13g2_fill_1 FILLER_41_155 ();
 sg13g2_fill_1 FILLER_41_164 ();
 sg13g2_fill_2 FILLER_41_188 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_fill_2 FILLER_41_223 ();
 sg13g2_fill_1 FILLER_41_225 ();
 sg13g2_fill_1 FILLER_41_247 ();
 sg13g2_fill_2 FILLER_41_253 ();
 sg13g2_decap_8 FILLER_41_291 ();
 sg13g2_decap_8 FILLER_41_298 ();
 sg13g2_fill_2 FILLER_41_305 ();
 sg13g2_fill_1 FILLER_41_307 ();
 sg13g2_decap_8 FILLER_41_313 ();
 sg13g2_decap_8 FILLER_41_320 ();
 sg13g2_decap_4 FILLER_41_339 ();
 sg13g2_fill_2 FILLER_41_343 ();
 sg13g2_decap_4 FILLER_41_351 ();
 sg13g2_decap_8 FILLER_41_367 ();
 sg13g2_decap_4 FILLER_41_405 ();
 sg13g2_decap_8 FILLER_42_0 ();
 sg13g2_fill_2 FILLER_42_7 ();
 sg13g2_fill_2 FILLER_42_22 ();
 sg13g2_fill_1 FILLER_42_24 ();
 sg13g2_fill_2 FILLER_42_33 ();
 sg13g2_decap_8 FILLER_42_47 ();
 sg13g2_fill_1 FILLER_42_54 ();
 sg13g2_fill_2 FILLER_42_68 ();
 sg13g2_fill_1 FILLER_42_70 ();
 sg13g2_fill_1 FILLER_42_109 ();
 sg13g2_fill_2 FILLER_42_120 ();
 sg13g2_fill_1 FILLER_42_122 ();
 sg13g2_fill_2 FILLER_42_139 ();
 sg13g2_decap_4 FILLER_42_147 ();
 sg13g2_fill_1 FILLER_42_151 ();
 sg13g2_fill_1 FILLER_42_181 ();
 sg13g2_decap_4 FILLER_42_202 ();
 sg13g2_fill_2 FILLER_42_206 ();
 sg13g2_decap_8 FILLER_42_226 ();
 sg13g2_fill_1 FILLER_42_233 ();
 sg13g2_decap_8 FILLER_42_239 ();
 sg13g2_fill_1 FILLER_42_246 ();
 sg13g2_decap_8 FILLER_42_251 ();
 sg13g2_fill_2 FILLER_42_258 ();
 sg13g2_fill_1 FILLER_42_260 ();
 sg13g2_decap_8 FILLER_42_282 ();
 sg13g2_decap_8 FILLER_42_289 ();
 sg13g2_decap_8 FILLER_42_296 ();
 sg13g2_fill_1 FILLER_42_303 ();
 sg13g2_fill_2 FILLER_42_320 ();
 sg13g2_fill_1 FILLER_42_322 ();
 sg13g2_decap_4 FILLER_42_329 ();
 sg13g2_fill_1 FILLER_42_338 ();
 sg13g2_fill_1 FILLER_42_345 ();
 sg13g2_fill_1 FILLER_42_352 ();
 sg13g2_decap_8 FILLER_42_371 ();
 sg13g2_fill_2 FILLER_42_378 ();
 sg13g2_fill_1 FILLER_42_385 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_4 FILLER_42_403 ();
 sg13g2_fill_2 FILLER_42_407 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_4 FILLER_43_7 ();
 sg13g2_fill_2 FILLER_43_11 ();
 sg13g2_decap_8 FILLER_43_17 ();
 sg13g2_fill_2 FILLER_43_24 ();
 sg13g2_fill_2 FILLER_43_30 ();
 sg13g2_fill_2 FILLER_43_57 ();
 sg13g2_decap_4 FILLER_43_71 ();
 sg13g2_fill_2 FILLER_43_75 ();
 sg13g2_decap_8 FILLER_43_101 ();
 sg13g2_decap_8 FILLER_43_108 ();
 sg13g2_fill_2 FILLER_43_115 ();
 sg13g2_decap_8 FILLER_43_139 ();
 sg13g2_decap_8 FILLER_43_146 ();
 sg13g2_fill_2 FILLER_43_153 ();
 sg13g2_fill_1 FILLER_43_155 ();
 sg13g2_decap_8 FILLER_43_200 ();
 sg13g2_decap_4 FILLER_43_207 ();
 sg13g2_fill_1 FILLER_43_216 ();
 sg13g2_fill_2 FILLER_43_227 ();
 sg13g2_fill_1 FILLER_43_229 ();
 sg13g2_fill_1 FILLER_43_260 ();
 sg13g2_fill_2 FILLER_43_265 ();
 sg13g2_fill_1 FILLER_43_267 ();
 sg13g2_decap_4 FILLER_43_274 ();
 sg13g2_fill_1 FILLER_43_278 ();
 sg13g2_fill_2 FILLER_43_284 ();
 sg13g2_fill_1 FILLER_43_286 ();
 sg13g2_fill_2 FILLER_43_302 ();
 sg13g2_fill_2 FILLER_43_309 ();
 sg13g2_fill_1 FILLER_43_311 ();
 sg13g2_decap_4 FILLER_43_317 ();
 sg13g2_fill_2 FILLER_43_321 ();
 sg13g2_decap_8 FILLER_43_327 ();
 sg13g2_decap_8 FILLER_43_334 ();
 sg13g2_decap_8 FILLER_43_341 ();
 sg13g2_decap_4 FILLER_43_348 ();
 sg13g2_fill_2 FILLER_43_352 ();
 sg13g2_decap_8 FILLER_43_368 ();
 sg13g2_decap_8 FILLER_43_375 ();
 sg13g2_decap_4 FILLER_43_382 ();
 sg13g2_fill_1 FILLER_43_386 ();
 sg13g2_fill_2 FILLER_43_391 ();
 sg13g2_decap_8 FILLER_43_398 ();
 sg13g2_decap_4 FILLER_43_405 ();
 sg13g2_fill_2 FILLER_44_0 ();
 sg13g2_fill_2 FILLER_44_12 ();
 sg13g2_fill_1 FILLER_44_14 ();
 sg13g2_decap_8 FILLER_44_31 ();
 sg13g2_decap_4 FILLER_44_41 ();
 sg13g2_decap_8 FILLER_44_50 ();
 sg13g2_decap_4 FILLER_44_79 ();
 sg13g2_fill_1 FILLER_44_83 ();
 sg13g2_decap_4 FILLER_44_103 ();
 sg13g2_fill_2 FILLER_44_107 ();
 sg13g2_decap_4 FILLER_44_117 ();
 sg13g2_fill_1 FILLER_44_121 ();
 sg13g2_decap_8 FILLER_44_136 ();
 sg13g2_decap_4 FILLER_44_143 ();
 sg13g2_decap_8 FILLER_44_153 ();
 sg13g2_fill_2 FILLER_44_160 ();
 sg13g2_fill_2 FILLER_44_182 ();
 sg13g2_fill_1 FILLER_44_184 ();
 sg13g2_fill_1 FILLER_44_195 ();
 sg13g2_decap_4 FILLER_44_202 ();
 sg13g2_decap_4 FILLER_44_224 ();
 sg13g2_fill_2 FILLER_44_245 ();
 sg13g2_fill_2 FILLER_44_271 ();
 sg13g2_decap_8 FILLER_44_286 ();
 sg13g2_fill_2 FILLER_44_309 ();
 sg13g2_fill_1 FILLER_44_311 ();
 sg13g2_fill_1 FILLER_44_324 ();
 sg13g2_fill_2 FILLER_44_331 ();
 sg13g2_fill_1 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_356 ();
 sg13g2_fill_1 FILLER_44_363 ();
 sg13g2_fill_2 FILLER_44_385 ();
 sg13g2_decap_8 FILLER_44_398 ();
 sg13g2_decap_4 FILLER_44_405 ();
 sg13g2_fill_1 FILLER_45_0 ();
 sg13g2_decap_4 FILLER_45_13 ();
 sg13g2_decap_8 FILLER_45_32 ();
 sg13g2_decap_4 FILLER_45_39 ();
 sg13g2_fill_2 FILLER_45_43 ();
 sg13g2_decap_4 FILLER_45_50 ();
 sg13g2_fill_2 FILLER_45_54 ();
 sg13g2_fill_2 FILLER_45_65 ();
 sg13g2_decap_8 FILLER_45_71 ();
 sg13g2_decap_8 FILLER_45_78 ();
 sg13g2_fill_2 FILLER_45_85 ();
 sg13g2_decap_8 FILLER_45_95 ();
 sg13g2_fill_2 FILLER_45_114 ();
 sg13g2_decap_8 FILLER_45_158 ();
 sg13g2_fill_1 FILLER_45_165 ();
 sg13g2_decap_8 FILLER_45_171 ();
 sg13g2_decap_8 FILLER_45_204 ();
 sg13g2_fill_2 FILLER_45_250 ();
 sg13g2_fill_1 FILLER_45_252 ();
 sg13g2_fill_2 FILLER_45_277 ();
 sg13g2_fill_2 FILLER_45_302 ();
 sg13g2_fill_1 FILLER_45_304 ();
 sg13g2_decap_4 FILLER_45_310 ();
 sg13g2_fill_2 FILLER_45_314 ();
 sg13g2_decap_8 FILLER_45_321 ();
 sg13g2_decap_8 FILLER_45_328 ();
 sg13g2_decap_8 FILLER_45_335 ();
 sg13g2_decap_8 FILLER_45_342 ();
 sg13g2_decap_4 FILLER_45_349 ();
 sg13g2_fill_2 FILLER_45_358 ();
 sg13g2_fill_1 FILLER_45_369 ();
 sg13g2_decap_8 FILLER_45_376 ();
 sg13g2_fill_1 FILLER_45_383 ();
 sg13g2_fill_2 FILLER_45_391 ();
 sg13g2_decap_4 FILLER_45_405 ();
 sg13g2_fill_1 FILLER_46_0 ();
 sg13g2_fill_2 FILLER_46_21 ();
 sg13g2_fill_1 FILLER_46_39 ();
 sg13g2_fill_2 FILLER_46_53 ();
 sg13g2_fill_1 FILLER_46_55 ();
 sg13g2_fill_1 FILLER_46_73 ();
 sg13g2_decap_4 FILLER_46_80 ();
 sg13g2_decap_4 FILLER_46_97 ();
 sg13g2_fill_2 FILLER_46_123 ();
 sg13g2_fill_1 FILLER_46_125 ();
 sg13g2_fill_1 FILLER_46_169 ();
 sg13g2_fill_2 FILLER_46_191 ();
 sg13g2_fill_1 FILLER_46_193 ();
 sg13g2_decap_8 FILLER_46_198 ();
 sg13g2_fill_1 FILLER_46_205 ();
 sg13g2_decap_4 FILLER_46_212 ();
 sg13g2_fill_1 FILLER_46_216 ();
 sg13g2_decap_4 FILLER_46_230 ();
 sg13g2_fill_2 FILLER_46_281 ();
 sg13g2_decap_8 FILLER_46_305 ();
 sg13g2_decap_8 FILLER_46_312 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_fill_2 FILLER_46_340 ();
 sg13g2_fill_1 FILLER_46_342 ();
 sg13g2_decap_4 FILLER_46_354 ();
 sg13g2_decap_4 FILLER_46_363 ();
 sg13g2_decap_8 FILLER_46_373 ();
 sg13g2_fill_2 FILLER_46_380 ();
 sg13g2_fill_2 FILLER_46_388 ();
 sg13g2_fill_1 FILLER_46_390 ();
 sg13g2_decap_8 FILLER_46_401 ();
 sg13g2_fill_1 FILLER_46_408 ();
 sg13g2_fill_1 FILLER_47_0 ();
 sg13g2_fill_1 FILLER_47_13 ();
 sg13g2_fill_1 FILLER_47_70 ();
 sg13g2_fill_2 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_127 ();
 sg13g2_decap_4 FILLER_47_134 ();
 sg13g2_fill_2 FILLER_47_173 ();
 sg13g2_fill_1 FILLER_47_175 ();
 sg13g2_fill_2 FILLER_47_184 ();
 sg13g2_fill_1 FILLER_47_186 ();
 sg13g2_fill_2 FILLER_47_191 ();
 sg13g2_fill_2 FILLER_47_202 ();
 sg13g2_decap_4 FILLER_47_208 ();
 sg13g2_decap_4 FILLER_47_228 ();
 sg13g2_fill_2 FILLER_47_300 ();
 sg13g2_fill_2 FILLER_47_314 ();
 sg13g2_fill_2 FILLER_47_322 ();
 sg13g2_fill_1 FILLER_47_324 ();
 sg13g2_fill_2 FILLER_47_335 ();
 sg13g2_fill_1 FILLER_47_337 ();
 sg13g2_decap_8 FILLER_47_349 ();
 sg13g2_decap_8 FILLER_47_356 ();
 sg13g2_decap_8 FILLER_47_363 ();
 sg13g2_decap_8 FILLER_47_376 ();
 sg13g2_decap_8 FILLER_47_383 ();
 sg13g2_decap_8 FILLER_47_390 ();
 sg13g2_fill_1 FILLER_47_397 ();
 sg13g2_decap_8 FILLER_47_402 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_12 ();
 sg13g2_fill_2 FILLER_48_19 ();
 sg13g2_fill_1 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_4 FILLER_48_49 ();
 sg13g2_fill_2 FILLER_48_73 ();
 sg13g2_fill_1 FILLER_48_75 ();
 sg13g2_fill_2 FILLER_48_112 ();
 sg13g2_fill_1 FILLER_48_114 ();
 sg13g2_decap_8 FILLER_48_120 ();
 sg13g2_decap_8 FILLER_48_127 ();
 sg13g2_decap_8 FILLER_48_134 ();
 sg13g2_decap_4 FILLER_48_141 ();
 sg13g2_fill_1 FILLER_48_145 ();
 sg13g2_decap_4 FILLER_48_163 ();
 sg13g2_fill_2 FILLER_48_181 ();
 sg13g2_fill_2 FILLER_48_191 ();
 sg13g2_fill_1 FILLER_48_193 ();
 sg13g2_fill_2 FILLER_48_203 ();
 sg13g2_fill_1 FILLER_48_205 ();
 sg13g2_fill_2 FILLER_48_270 ();
 sg13g2_fill_1 FILLER_48_278 ();
 sg13g2_fill_2 FILLER_48_307 ();
 sg13g2_decap_4 FILLER_48_314 ();
 sg13g2_fill_1 FILLER_48_318 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_4 FILLER_48_350 ();
 sg13g2_fill_1 FILLER_48_354 ();
 sg13g2_decap_8 FILLER_48_359 ();
 sg13g2_fill_2 FILLER_48_366 ();
 sg13g2_fill_2 FILLER_48_378 ();
 sg13g2_fill_1 FILLER_48_380 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_fill_2 FILLER_48_406 ();
 sg13g2_fill_1 FILLER_48_408 ();
 sg13g2_decap_4 FILLER_49_0 ();
 sg13g2_fill_1 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_fill_2 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_fill_2 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_77 ();
 sg13g2_decap_8 FILLER_49_97 ();
 sg13g2_decap_4 FILLER_49_104 ();
 sg13g2_fill_1 FILLER_49_108 ();
 sg13g2_decap_4 FILLER_49_129 ();
 sg13g2_fill_2 FILLER_49_133 ();
 sg13g2_decap_8 FILLER_49_141 ();
 sg13g2_decap_4 FILLER_49_148 ();
 sg13g2_fill_1 FILLER_49_152 ();
 sg13g2_decap_4 FILLER_49_169 ();
 sg13g2_fill_1 FILLER_49_173 ();
 sg13g2_decap_4 FILLER_49_178 ();
 sg13g2_fill_1 FILLER_49_182 ();
 sg13g2_decap_4 FILLER_49_188 ();
 sg13g2_decap_4 FILLER_49_207 ();
 sg13g2_fill_1 FILLER_49_211 ();
 sg13g2_fill_2 FILLER_49_220 ();
 sg13g2_fill_2 FILLER_49_234 ();
 sg13g2_fill_1 FILLER_49_262 ();
 sg13g2_decap_4 FILLER_49_276 ();
 sg13g2_fill_1 FILLER_49_280 ();
 sg13g2_decap_4 FILLER_49_307 ();
 sg13g2_fill_2 FILLER_49_319 ();
 sg13g2_decap_4 FILLER_49_326 ();
 sg13g2_fill_1 FILLER_49_334 ();
 sg13g2_fill_1 FILLER_49_347 ();
 sg13g2_decap_4 FILLER_49_376 ();
 sg13g2_fill_2 FILLER_49_380 ();
 sg13g2_decap_4 FILLER_49_391 ();
 sg13g2_decap_8 FILLER_49_400 ();
 sg13g2_fill_2 FILLER_49_407 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_fill_1 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_13 ();
 sg13g2_fill_2 FILLER_50_33 ();
 sg13g2_fill_1 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_53 ();
 sg13g2_fill_2 FILLER_50_60 ();
 sg13g2_fill_1 FILLER_50_62 ();
 sg13g2_decap_8 FILLER_50_75 ();
 sg13g2_fill_2 FILLER_50_82 ();
 sg13g2_decap_8 FILLER_50_101 ();
 sg13g2_fill_2 FILLER_50_136 ();
 sg13g2_fill_1 FILLER_50_138 ();
 sg13g2_decap_4 FILLER_50_149 ();
 sg13g2_fill_1 FILLER_50_153 ();
 sg13g2_decap_8 FILLER_50_159 ();
 sg13g2_fill_2 FILLER_50_166 ();
 sg13g2_decap_8 FILLER_50_177 ();
 sg13g2_fill_2 FILLER_50_184 ();
 sg13g2_decap_8 FILLER_50_191 ();
 sg13g2_decap_8 FILLER_50_198 ();
 sg13g2_fill_1 FILLER_50_205 ();
 sg13g2_fill_2 FILLER_50_212 ();
 sg13g2_fill_1 FILLER_50_214 ();
 sg13g2_decap_8 FILLER_50_225 ();
 sg13g2_fill_1 FILLER_50_232 ();
 sg13g2_fill_2 FILLER_50_255 ();
 sg13g2_fill_1 FILLER_50_257 ();
 sg13g2_decap_4 FILLER_50_276 ();
 sg13g2_fill_1 FILLER_50_280 ();
 sg13g2_fill_2 FILLER_50_292 ();
 sg13g2_fill_1 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_318 ();
 sg13g2_decap_8 FILLER_50_325 ();
 sg13g2_fill_2 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_351 ();
 sg13g2_fill_2 FILLER_50_358 ();
 sg13g2_fill_1 FILLER_50_360 ();
 sg13g2_decap_8 FILLER_50_369 ();
 sg13g2_decap_8 FILLER_50_376 ();
 sg13g2_decap_8 FILLER_50_383 ();
 sg13g2_decap_8 FILLER_50_390 ();
 sg13g2_decap_8 FILLER_50_397 ();
 sg13g2_decap_4 FILLER_50_404 ();
 sg13g2_fill_1 FILLER_50_408 ();
 sg13g2_decap_4 FILLER_51_13 ();
 sg13g2_fill_2 FILLER_51_30 ();
 sg13g2_fill_1 FILLER_51_32 ();
 sg13g2_fill_2 FILLER_51_99 ();
 sg13g2_fill_1 FILLER_51_101 ();
 sg13g2_fill_1 FILLER_51_139 ();
 sg13g2_fill_2 FILLER_51_157 ();
 sg13g2_decap_8 FILLER_51_169 ();
 sg13g2_fill_2 FILLER_51_176 ();
 sg13g2_fill_1 FILLER_51_178 ();
 sg13g2_fill_2 FILLER_51_183 ();
 sg13g2_fill_2 FILLER_51_201 ();
 sg13g2_fill_2 FILLER_51_216 ();
 sg13g2_decap_8 FILLER_51_223 ();
 sg13g2_fill_2 FILLER_51_230 ();
 sg13g2_fill_1 FILLER_51_232 ();
 sg13g2_fill_1 FILLER_51_237 ();
 sg13g2_decap_4 FILLER_51_252 ();
 sg13g2_fill_1 FILLER_51_256 ();
 sg13g2_decap_4 FILLER_51_262 ();
 sg13g2_decap_4 FILLER_51_275 ();
 sg13g2_decap_8 FILLER_51_283 ();
 sg13g2_decap_8 FILLER_51_290 ();
 sg13g2_fill_2 FILLER_51_297 ();
 sg13g2_fill_1 FILLER_51_299 ();
 sg13g2_decap_8 FILLER_51_309 ();
 sg13g2_decap_4 FILLER_51_316 ();
 sg13g2_fill_2 FILLER_51_320 ();
 sg13g2_fill_2 FILLER_51_333 ();
 sg13g2_decap_8 FILLER_51_346 ();
 sg13g2_fill_2 FILLER_51_353 ();
 sg13g2_fill_1 FILLER_51_355 ();
 sg13g2_fill_2 FILLER_51_365 ();
 sg13g2_fill_1 FILLER_51_367 ();
 sg13g2_decap_8 FILLER_51_374 ();
 sg13g2_fill_2 FILLER_51_381 ();
 sg13g2_fill_1 FILLER_51_383 ();
 sg13g2_decap_8 FILLER_51_401 ();
 sg13g2_fill_1 FILLER_51_408 ();
 sg13g2_fill_1 FILLER_52_0 ();
 sg13g2_fill_1 FILLER_52_16 ();
 sg13g2_decap_8 FILLER_52_25 ();
 sg13g2_decap_4 FILLER_52_32 ();
 sg13g2_fill_1 FILLER_52_36 ();
 sg13g2_fill_1 FILLER_52_45 ();
 sg13g2_decap_8 FILLER_52_54 ();
 sg13g2_fill_1 FILLER_52_61 ();
 sg13g2_fill_2 FILLER_52_83 ();
 sg13g2_fill_1 FILLER_52_94 ();
 sg13g2_fill_1 FILLER_52_103 ();
 sg13g2_decap_8 FILLER_52_109 ();
 sg13g2_fill_2 FILLER_52_116 ();
 sg13g2_fill_1 FILLER_52_118 ();
 sg13g2_fill_1 FILLER_52_164 ();
 sg13g2_fill_1 FILLER_52_197 ();
 sg13g2_decap_4 FILLER_52_212 ();
 sg13g2_fill_1 FILLER_52_216 ();
 sg13g2_fill_2 FILLER_52_249 ();
 sg13g2_fill_1 FILLER_52_251 ();
 sg13g2_fill_2 FILLER_52_270 ();
 sg13g2_fill_2 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_309 ();
 sg13g2_decap_4 FILLER_52_316 ();
 sg13g2_fill_1 FILLER_52_320 ();
 sg13g2_fill_1 FILLER_52_326 ();
 sg13g2_decap_8 FILLER_52_331 ();
 sg13g2_decap_8 FILLER_52_338 ();
 sg13g2_decap_4 FILLER_52_345 ();
 sg13g2_fill_2 FILLER_52_349 ();
 sg13g2_fill_2 FILLER_52_371 ();
 sg13g2_fill_1 FILLER_52_373 ();
 sg13g2_decap_8 FILLER_52_379 ();
 sg13g2_fill_1 FILLER_52_386 ();
 sg13g2_decap_8 FILLER_52_398 ();
 sg13g2_decap_4 FILLER_52_405 ();
 sg13g2_fill_2 FILLER_53_0 ();
 sg13g2_fill_2 FILLER_53_14 ();
 sg13g2_fill_1 FILLER_53_33 ();
 sg13g2_decap_4 FILLER_53_42 ();
 sg13g2_fill_1 FILLER_53_46 ();
 sg13g2_decap_8 FILLER_53_59 ();
 sg13g2_decap_4 FILLER_53_66 ();
 sg13g2_fill_2 FILLER_53_93 ();
 sg13g2_fill_2 FILLER_53_100 ();
 sg13g2_decap_8 FILLER_53_111 ();
 sg13g2_decap_4 FILLER_53_118 ();
 sg13g2_fill_2 FILLER_53_122 ();
 sg13g2_fill_2 FILLER_53_128 ();
 sg13g2_fill_2 FILLER_53_134 ();
 sg13g2_decap_4 FILLER_53_178 ();
 sg13g2_fill_2 FILLER_53_182 ();
 sg13g2_fill_2 FILLER_53_189 ();
 sg13g2_fill_1 FILLER_53_191 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_4 FILLER_53_217 ();
 sg13g2_fill_1 FILLER_53_238 ();
 sg13g2_fill_1 FILLER_53_252 ();
 sg13g2_fill_1 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_286 ();
 sg13g2_decap_4 FILLER_53_293 ();
 sg13g2_fill_1 FILLER_53_301 ();
 sg13g2_fill_2 FILLER_53_307 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_fill_2 FILLER_53_322 ();
 sg13g2_fill_1 FILLER_53_324 ();
 sg13g2_decap_4 FILLER_53_338 ();
 sg13g2_fill_2 FILLER_53_342 ();
 sg13g2_decap_8 FILLER_53_349 ();
 sg13g2_decap_8 FILLER_53_356 ();
 sg13g2_decap_4 FILLER_53_363 ();
 sg13g2_fill_1 FILLER_53_367 ();
 sg13g2_decap_8 FILLER_53_376 ();
 sg13g2_decap_8 FILLER_53_383 ();
 sg13g2_fill_2 FILLER_53_390 ();
 sg13g2_decap_8 FILLER_53_396 ();
 sg13g2_decap_4 FILLER_53_403 ();
 sg13g2_fill_2 FILLER_53_407 ();
 sg13g2_decap_8 FILLER_54_0 ();
 sg13g2_fill_1 FILLER_54_7 ();
 sg13g2_fill_2 FILLER_54_15 ();
 sg13g2_decap_4 FILLER_54_30 ();
 sg13g2_decap_4 FILLER_54_42 ();
 sg13g2_fill_2 FILLER_54_51 ();
 sg13g2_fill_1 FILLER_54_53 ();
 sg13g2_decap_8 FILLER_54_62 ();
 sg13g2_decap_8 FILLER_54_69 ();
 sg13g2_decap_8 FILLER_54_76 ();
 sg13g2_decap_4 FILLER_54_118 ();
 sg13g2_fill_1 FILLER_54_122 ();
 sg13g2_decap_4 FILLER_54_137 ();
 sg13g2_fill_2 FILLER_54_147 ();
 sg13g2_fill_1 FILLER_54_149 ();
 sg13g2_fill_1 FILLER_54_158 ();
 sg13g2_decap_8 FILLER_54_169 ();
 sg13g2_decap_8 FILLER_54_176 ();
 sg13g2_decap_8 FILLER_54_183 ();
 sg13g2_decap_4 FILLER_54_190 ();
 sg13g2_fill_1 FILLER_54_194 ();
 sg13g2_decap_8 FILLER_54_206 ();
 sg13g2_decap_8 FILLER_54_213 ();
 sg13g2_decap_4 FILLER_54_220 ();
 sg13g2_fill_2 FILLER_54_224 ();
 sg13g2_decap_8 FILLER_54_286 ();
 sg13g2_fill_2 FILLER_54_293 ();
 sg13g2_fill_1 FILLER_54_295 ();
 sg13g2_decap_8 FILLER_54_302 ();
 sg13g2_decap_8 FILLER_54_309 ();
 sg13g2_fill_1 FILLER_54_316 ();
 sg13g2_decap_8 FILLER_54_324 ();
 sg13g2_fill_2 FILLER_54_331 ();
 sg13g2_fill_1 FILLER_54_333 ();
 sg13g2_decap_8 FILLER_54_344 ();
 sg13g2_decap_8 FILLER_54_351 ();
 sg13g2_decap_8 FILLER_54_358 ();
 sg13g2_decap_8 FILLER_54_365 ();
 sg13g2_decap_8 FILLER_54_377 ();
 sg13g2_fill_1 FILLER_55_0 ();
 sg13g2_decap_4 FILLER_55_12 ();
 sg13g2_fill_2 FILLER_55_43 ();
 sg13g2_decap_8 FILLER_55_66 ();
 sg13g2_decap_8 FILLER_55_73 ();
 sg13g2_decap_4 FILLER_55_80 ();
 sg13g2_fill_1 FILLER_55_106 ();
 sg13g2_fill_2 FILLER_55_118 ();
 sg13g2_fill_1 FILLER_55_120 ();
 sg13g2_fill_1 FILLER_55_142 ();
 sg13g2_decap_8 FILLER_55_151 ();
 sg13g2_decap_8 FILLER_55_158 ();
 sg13g2_fill_1 FILLER_55_165 ();
 sg13g2_decap_4 FILLER_55_183 ();
 sg13g2_fill_2 FILLER_55_187 ();
 sg13g2_decap_8 FILLER_55_214 ();
 sg13g2_decap_8 FILLER_55_221 ();
 sg13g2_fill_1 FILLER_55_254 ();
 sg13g2_fill_1 FILLER_55_262 ();
 sg13g2_fill_2 FILLER_55_283 ();
 sg13g2_fill_1 FILLER_55_285 ();
 sg13g2_fill_1 FILLER_55_305 ();
 sg13g2_fill_2 FILLER_55_316 ();
 sg13g2_fill_2 FILLER_55_373 ();
 sg13g2_fill_1 FILLER_55_375 ();
 sg13g2_decap_8 FILLER_55_382 ();
 sg13g2_decap_8 FILLER_55_389 ();
 sg13g2_decap_8 FILLER_55_401 ();
 sg13g2_fill_1 FILLER_55_408 ();
 sg13g2_fill_1 FILLER_56_0 ();
 sg13g2_decap_4 FILLER_56_13 ();
 sg13g2_fill_1 FILLER_56_46 ();
 sg13g2_fill_1 FILLER_56_54 ();
 sg13g2_fill_2 FILLER_56_65 ();
 sg13g2_fill_1 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_79 ();
 sg13g2_fill_2 FILLER_56_86 ();
 sg13g2_fill_1 FILLER_56_88 ();
 sg13g2_decap_4 FILLER_56_102 ();
 sg13g2_fill_2 FILLER_56_114 ();
 sg13g2_decap_8 FILLER_56_146 ();
 sg13g2_fill_2 FILLER_56_153 ();
 sg13g2_decap_4 FILLER_56_166 ();
 sg13g2_decap_8 FILLER_56_223 ();
 sg13g2_fill_1 FILLER_56_230 ();
 sg13g2_fill_1 FILLER_56_271 ();
 sg13g2_fill_2 FILLER_56_279 ();
 sg13g2_fill_1 FILLER_56_281 ();
 sg13g2_fill_1 FILLER_56_306 ();
 sg13g2_decap_4 FILLER_56_326 ();
 sg13g2_fill_2 FILLER_56_330 ();
 sg13g2_fill_1 FILLER_56_344 ();
 sg13g2_fill_2 FILLER_56_353 ();
 sg13g2_decap_8 FILLER_56_361 ();
 sg13g2_decap_8 FILLER_56_368 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_fill_2 FILLER_56_406 ();
 sg13g2_fill_1 FILLER_56_408 ();
 sg13g2_fill_2 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_29 ();
 sg13g2_fill_1 FILLER_57_36 ();
 sg13g2_fill_2 FILLER_57_89 ();
 sg13g2_fill_1 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_100 ();
 sg13g2_decap_8 FILLER_57_115 ();
 sg13g2_fill_2 FILLER_57_122 ();
 sg13g2_fill_1 FILLER_57_139 ();
 sg13g2_fill_2 FILLER_57_150 ();
 sg13g2_fill_1 FILLER_57_152 ();
 sg13g2_fill_1 FILLER_57_163 ();
 sg13g2_decap_4 FILLER_57_191 ();
 sg13g2_fill_2 FILLER_57_200 ();
 sg13g2_fill_1 FILLER_57_202 ();
 sg13g2_fill_1 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_226 ();
 sg13g2_decap_8 FILLER_57_233 ();
 sg13g2_decap_8 FILLER_57_240 ();
 sg13g2_decap_4 FILLER_57_247 ();
 sg13g2_fill_2 FILLER_57_251 ();
 sg13g2_fill_2 FILLER_57_283 ();
 sg13g2_decap_8 FILLER_57_293 ();
 sg13g2_decap_4 FILLER_57_305 ();
 sg13g2_fill_1 FILLER_57_313 ();
 sg13g2_decap_8 FILLER_57_319 ();
 sg13g2_decap_8 FILLER_57_326 ();
 sg13g2_decap_8 FILLER_57_333 ();
 sg13g2_fill_1 FILLER_57_340 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_fill_1 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_370 ();
 sg13g2_fill_2 FILLER_57_377 ();
 sg13g2_decap_8 FILLER_57_388 ();
 sg13g2_decap_8 FILLER_57_395 ();
 sg13g2_decap_8 FILLER_57_402 ();
 sg13g2_fill_1 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_22 ();
 sg13g2_decap_8 FILLER_58_29 ();
 sg13g2_decap_8 FILLER_58_36 ();
 sg13g2_fill_2 FILLER_58_43 ();
 sg13g2_fill_1 FILLER_58_45 ();
 sg13g2_decap_4 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_65 ();
 sg13g2_fill_2 FILLER_58_72 ();
 sg13g2_decap_8 FILLER_58_108 ();
 sg13g2_decap_4 FILLER_58_115 ();
 sg13g2_fill_2 FILLER_58_138 ();
 sg13g2_fill_1 FILLER_58_140 ();
 sg13g2_fill_2 FILLER_58_166 ();
 sg13g2_decap_8 FILLER_58_186 ();
 sg13g2_decap_4 FILLER_58_193 ();
 sg13g2_fill_2 FILLER_58_197 ();
 sg13g2_decap_8 FILLER_58_235 ();
 sg13g2_fill_2 FILLER_58_242 ();
 sg13g2_fill_1 FILLER_58_244 ();
 sg13g2_fill_2 FILLER_58_272 ();
 sg13g2_fill_1 FILLER_58_274 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_fill_1 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_342 ();
 sg13g2_decap_8 FILLER_58_349 ();
 sg13g2_decap_8 FILLER_58_356 ();
 sg13g2_fill_2 FILLER_58_363 ();
 sg13g2_fill_1 FILLER_58_365 ();
 sg13g2_decap_8 FILLER_58_370 ();
 sg13g2_decap_8 FILLER_58_377 ();
 sg13g2_decap_8 FILLER_58_384 ();
 sg13g2_fill_1 FILLER_58_391 ();
 sg13g2_decap_8 FILLER_58_397 ();
 sg13g2_decap_4 FILLER_58_404 ();
 sg13g2_fill_1 FILLER_58_408 ();
 sg13g2_decap_4 FILLER_59_0 ();
 sg13g2_fill_1 FILLER_59_4 ();
 sg13g2_decap_8 FILLER_59_15 ();
 sg13g2_decap_8 FILLER_59_22 ();
 sg13g2_decap_8 FILLER_59_29 ();
 sg13g2_decap_8 FILLER_59_36 ();
 sg13g2_decap_8 FILLER_59_43 ();
 sg13g2_decap_8 FILLER_59_50 ();
 sg13g2_decap_8 FILLER_59_57 ();
 sg13g2_decap_8 FILLER_59_64 ();
 sg13g2_decap_8 FILLER_59_71 ();
 sg13g2_fill_2 FILLER_59_78 ();
 sg13g2_decap_4 FILLER_59_86 ();
 sg13g2_fill_1 FILLER_59_103 ();
 sg13g2_fill_2 FILLER_59_117 ();
 sg13g2_fill_2 FILLER_59_137 ();
 sg13g2_fill_1 FILLER_59_139 ();
 sg13g2_fill_1 FILLER_59_148 ();
 sg13g2_decap_4 FILLER_59_163 ();
 sg13g2_fill_1 FILLER_59_167 ();
 sg13g2_decap_8 FILLER_59_177 ();
 sg13g2_decap_8 FILLER_59_184 ();
 sg13g2_decap_8 FILLER_59_191 ();
 sg13g2_fill_2 FILLER_59_198 ();
 sg13g2_fill_2 FILLER_59_217 ();
 sg13g2_decap_8 FILLER_59_241 ();
 sg13g2_fill_2 FILLER_59_265 ();
 sg13g2_decap_8 FILLER_59_272 ();
 sg13g2_fill_2 FILLER_59_279 ();
 sg13g2_fill_1 FILLER_59_281 ();
 sg13g2_fill_2 FILLER_59_290 ();
 sg13g2_fill_2 FILLER_59_314 ();
 sg13g2_decap_4 FILLER_59_320 ();
 sg13g2_fill_2 FILLER_59_324 ();
 sg13g2_fill_1 FILLER_59_342 ();
 sg13g2_decap_4 FILLER_59_351 ();
 sg13g2_fill_2 FILLER_59_360 ();
 sg13g2_fill_1 FILLER_59_362 ();
 sg13g2_fill_2 FILLER_59_368 ();
 sg13g2_fill_1 FILLER_59_370 ();
 sg13g2_fill_1 FILLER_59_378 ();
 sg13g2_fill_1 FILLER_59_408 ();
 sg13g2_decap_4 FILLER_60_0 ();
 sg13g2_decap_4 FILLER_60_24 ();
 sg13g2_fill_2 FILLER_60_28 ();
 sg13g2_fill_2 FILLER_60_48 ();
 sg13g2_decap_8 FILLER_60_55 ();
 sg13g2_decap_4 FILLER_60_62 ();
 sg13g2_fill_2 FILLER_60_66 ();
 sg13g2_decap_8 FILLER_60_111 ();
 sg13g2_fill_1 FILLER_60_155 ();
 sg13g2_fill_2 FILLER_60_160 ();
 sg13g2_fill_1 FILLER_60_162 ();
 sg13g2_fill_1 FILLER_60_174 ();
 sg13g2_fill_2 FILLER_60_197 ();
 sg13g2_decap_4 FILLER_60_214 ();
 sg13g2_fill_1 FILLER_60_227 ();
 sg13g2_fill_2 FILLER_60_281 ();
 sg13g2_fill_1 FILLER_60_283 ();
 sg13g2_decap_8 FILLER_60_345 ();
 sg13g2_decap_4 FILLER_60_352 ();
 sg13g2_fill_1 FILLER_60_356 ();
 sg13g2_fill_2 FILLER_60_374 ();
 sg13g2_fill_1 FILLER_60_376 ();
 sg13g2_decap_4 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_398 ();
 sg13g2_decap_4 FILLER_60_405 ();
 sg13g2_fill_1 FILLER_61_0 ();
 sg13g2_fill_1 FILLER_61_18 ();
 sg13g2_fill_1 FILLER_61_39 ();
 sg13g2_fill_2 FILLER_61_55 ();
 sg13g2_fill_1 FILLER_61_57 ();
 sg13g2_decap_8 FILLER_61_70 ();
 sg13g2_fill_2 FILLER_61_77 ();
 sg13g2_fill_1 FILLER_61_79 ();
 sg13g2_decap_8 FILLER_61_91 ();
 sg13g2_fill_1 FILLER_61_103 ();
 sg13g2_decap_8 FILLER_61_109 ();
 sg13g2_decap_4 FILLER_61_116 ();
 sg13g2_fill_2 FILLER_61_120 ();
 sg13g2_decap_4 FILLER_61_173 ();
 sg13g2_fill_1 FILLER_61_185 ();
 sg13g2_fill_1 FILLER_61_204 ();
 sg13g2_decap_4 FILLER_61_209 ();
 sg13g2_fill_1 FILLER_61_213 ();
 sg13g2_fill_2 FILLER_61_222 ();
 sg13g2_fill_1 FILLER_61_224 ();
 sg13g2_fill_1 FILLER_61_235 ();
 sg13g2_fill_1 FILLER_61_271 ();
 sg13g2_decap_4 FILLER_61_281 ();
 sg13g2_fill_2 FILLER_61_291 ();
 sg13g2_fill_1 FILLER_61_293 ();
 sg13g2_fill_2 FILLER_61_330 ();
 sg13g2_fill_1 FILLER_61_337 ();
 sg13g2_fill_1 FILLER_61_354 ();
 sg13g2_decap_4 FILLER_61_370 ();
 sg13g2_decap_4 FILLER_61_386 ();
 sg13g2_decap_8 FILLER_61_401 ();
 sg13g2_fill_1 FILLER_61_408 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_fill_2 FILLER_62_23 ();
 sg13g2_fill_2 FILLER_62_57 ();
 sg13g2_decap_8 FILLER_62_80 ();
 sg13g2_decap_8 FILLER_62_87 ();
 sg13g2_fill_2 FILLER_62_94 ();
 sg13g2_fill_2 FILLER_62_108 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_fill_1 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_143 ();
 sg13g2_decap_4 FILLER_62_150 ();
 sg13g2_fill_2 FILLER_62_154 ();
 sg13g2_fill_1 FILLER_62_164 ();
 sg13g2_fill_1 FILLER_62_169 ();
 sg13g2_fill_2 FILLER_62_180 ();
 sg13g2_fill_2 FILLER_62_199 ();
 sg13g2_fill_1 FILLER_62_205 ();
 sg13g2_fill_1 FILLER_62_218 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_4 FILLER_62_231 ();
 sg13g2_fill_1 FILLER_62_235 ();
 sg13g2_fill_1 FILLER_62_283 ();
 sg13g2_fill_2 FILLER_62_300 ();
 sg13g2_fill_1 FILLER_62_302 ();
 sg13g2_fill_2 FILLER_62_311 ();
 sg13g2_fill_1 FILLER_62_313 ();
 sg13g2_fill_2 FILLER_62_325 ();
 sg13g2_fill_1 FILLER_62_327 ();
 sg13g2_fill_1 FILLER_62_333 ();
 sg13g2_fill_1 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_361 ();
 sg13g2_fill_1 FILLER_62_368 ();
 sg13g2_decap_8 FILLER_62_374 ();
 sg13g2_decap_8 FILLER_62_381 ();
 sg13g2_decap_8 FILLER_62_388 ();
 sg13g2_fill_2 FILLER_62_406 ();
 sg13g2_fill_1 FILLER_62_408 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_fill_2 FILLER_63_7 ();
 sg13g2_fill_1 FILLER_63_9 ();
 sg13g2_fill_1 FILLER_63_34 ();
 sg13g2_fill_1 FILLER_63_44 ();
 sg13g2_fill_2 FILLER_63_49 ();
 sg13g2_fill_1 FILLER_63_51 ();
 sg13g2_decap_4 FILLER_63_77 ();
 sg13g2_fill_2 FILLER_63_87 ();
 sg13g2_fill_1 FILLER_63_89 ();
 sg13g2_fill_1 FILLER_63_110 ();
 sg13g2_fill_1 FILLER_63_135 ();
 sg13g2_fill_1 FILLER_63_146 ();
 sg13g2_decap_8 FILLER_63_155 ();
 sg13g2_decap_8 FILLER_63_162 ();
 sg13g2_decap_8 FILLER_63_169 ();
 sg13g2_decap_8 FILLER_63_176 ();
 sg13g2_fill_2 FILLER_63_183 ();
 sg13g2_fill_2 FILLER_63_191 ();
 sg13g2_fill_1 FILLER_63_193 ();
 sg13g2_fill_2 FILLER_63_199 ();
 sg13g2_fill_1 FILLER_63_201 ();
 sg13g2_fill_2 FILLER_63_206 ();
 sg13g2_fill_1 FILLER_63_208 ();
 sg13g2_decap_8 FILLER_63_232 ();
 sg13g2_decap_4 FILLER_63_239 ();
 sg13g2_fill_2 FILLER_63_243 ();
 sg13g2_fill_1 FILLER_63_253 ();
 sg13g2_decap_8 FILLER_63_264 ();
 sg13g2_decap_4 FILLER_63_276 ();
 sg13g2_fill_2 FILLER_63_293 ();
 sg13g2_fill_1 FILLER_63_295 ();
 sg13g2_decap_4 FILLER_63_309 ();
 sg13g2_decap_8 FILLER_63_319 ();
 sg13g2_decap_4 FILLER_63_326 ();
 sg13g2_fill_1 FILLER_63_330 ();
 sg13g2_fill_2 FILLER_63_349 ();
 sg13g2_decap_8 FILLER_63_355 ();
 sg13g2_decap_8 FILLER_63_362 ();
 sg13g2_decap_4 FILLER_63_369 ();
 sg13g2_fill_1 FILLER_63_373 ();
 sg13g2_decap_4 FILLER_63_379 ();
 sg13g2_decap_8 FILLER_63_388 ();
 sg13g2_decap_8 FILLER_63_395 ();
 sg13g2_decap_8 FILLER_63_402 ();
 sg13g2_decap_8 FILLER_64_0 ();
 sg13g2_decap_8 FILLER_64_7 ();
 sg13g2_decap_4 FILLER_64_14 ();
 sg13g2_decap_8 FILLER_64_34 ();
 sg13g2_decap_8 FILLER_64_41 ();
 sg13g2_decap_8 FILLER_64_74 ();
 sg13g2_fill_1 FILLER_64_81 ();
 sg13g2_decap_4 FILLER_64_93 ();
 sg13g2_fill_2 FILLER_64_97 ();
 sg13g2_fill_1 FILLER_64_116 ();
 sg13g2_decap_4 FILLER_64_160 ();
 sg13g2_fill_2 FILLER_64_183 ();
 sg13g2_fill_1 FILLER_64_185 ();
 sg13g2_fill_2 FILLER_64_198 ();
 sg13g2_fill_1 FILLER_64_200 ();
 sg13g2_fill_1 FILLER_64_218 ();
 sg13g2_decap_8 FILLER_64_239 ();
 sg13g2_decap_8 FILLER_64_246 ();
 sg13g2_fill_1 FILLER_64_253 ();
 sg13g2_decap_4 FILLER_64_268 ();
 sg13g2_fill_2 FILLER_64_284 ();
 sg13g2_decap_4 FILLER_64_290 ();
 sg13g2_fill_1 FILLER_64_294 ();
 sg13g2_decap_8 FILLER_64_300 ();
 sg13g2_decap_8 FILLER_64_307 ();
 sg13g2_decap_4 FILLER_64_314 ();
 sg13g2_fill_1 FILLER_64_318 ();
 sg13g2_decap_8 FILLER_64_332 ();
 sg13g2_fill_2 FILLER_64_339 ();
 sg13g2_fill_1 FILLER_64_341 ();
 sg13g2_fill_2 FILLER_64_346 ();
 sg13g2_fill_2 FILLER_64_359 ();
 sg13g2_fill_1 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_4 FILLER_64_403 ();
 sg13g2_fill_2 FILLER_64_407 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_fill_2 FILLER_65_27 ();
 sg13g2_decap_8 FILLER_65_47 ();
 sg13g2_fill_1 FILLER_65_62 ();
 sg13g2_decap_8 FILLER_65_68 ();
 sg13g2_decap_4 FILLER_65_75 ();
 sg13g2_fill_1 FILLER_65_79 ();
 sg13g2_decap_8 FILLER_65_92 ();
 sg13g2_decap_4 FILLER_65_99 ();
 sg13g2_fill_1 FILLER_65_103 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_fill_1 FILLER_65_126 ();
 sg13g2_fill_1 FILLER_65_154 ();
 sg13g2_fill_2 FILLER_65_201 ();
 sg13g2_fill_2 FILLER_65_215 ();
 sg13g2_fill_1 FILLER_65_247 ();
 sg13g2_fill_1 FILLER_65_253 ();
 sg13g2_decap_8 FILLER_65_274 ();
 sg13g2_decap_8 FILLER_65_281 ();
 sg13g2_fill_1 FILLER_65_288 ();
 sg13g2_fill_2 FILLER_65_293 ();
 sg13g2_fill_1 FILLER_65_307 ();
 sg13g2_fill_1 FILLER_65_313 ();
 sg13g2_decap_8 FILLER_65_319 ();
 sg13g2_decap_8 FILLER_65_326 ();
 sg13g2_decap_8 FILLER_65_333 ();
 sg13g2_fill_2 FILLER_65_340 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_fill_2 FILLER_65_357 ();
 sg13g2_fill_1 FILLER_65_391 ();
 sg13g2_fill_2 FILLER_65_406 ();
 sg13g2_fill_1 FILLER_65_408 ();
 sg13g2_decap_8 FILLER_66_0 ();
 sg13g2_decap_8 FILLER_66_7 ();
 sg13g2_fill_2 FILLER_66_14 ();
 sg13g2_fill_1 FILLER_66_16 ();
 sg13g2_decap_8 FILLER_66_22 ();
 sg13g2_decap_8 FILLER_66_29 ();
 sg13g2_decap_8 FILLER_66_36 ();
 sg13g2_decap_8 FILLER_66_43 ();
 sg13g2_fill_1 FILLER_66_50 ();
 sg13g2_decap_4 FILLER_66_55 ();
 sg13g2_fill_2 FILLER_66_59 ();
 sg13g2_decap_4 FILLER_66_66 ();
 sg13g2_fill_2 FILLER_66_70 ();
 sg13g2_fill_2 FILLER_66_93 ();
 sg13g2_fill_1 FILLER_66_95 ();
 sg13g2_decap_8 FILLER_66_109 ();
 sg13g2_decap_4 FILLER_66_116 ();
 sg13g2_decap_8 FILLER_66_128 ();
 sg13g2_fill_2 FILLER_66_135 ();
 sg13g2_fill_1 FILLER_66_137 ();
 sg13g2_fill_2 FILLER_66_143 ();
 sg13g2_fill_1 FILLER_66_145 ();
 sg13g2_fill_2 FILLER_66_177 ();
 sg13g2_fill_2 FILLER_66_187 ();
 sg13g2_decap_4 FILLER_66_219 ();
 sg13g2_fill_1 FILLER_66_223 ();
 sg13g2_decap_8 FILLER_66_230 ();
 sg13g2_fill_1 FILLER_66_237 ();
 sg13g2_decap_8 FILLER_66_261 ();
 sg13g2_decap_4 FILLER_66_268 ();
 sg13g2_fill_1 FILLER_66_272 ();
 sg13g2_fill_1 FILLER_66_286 ();
 sg13g2_decap_4 FILLER_66_296 ();
 sg13g2_fill_2 FILLER_66_306 ();
 sg13g2_decap_8 FILLER_66_336 ();
 sg13g2_decap_4 FILLER_66_343 ();
 sg13g2_fill_1 FILLER_66_347 ();
 sg13g2_fill_2 FILLER_66_354 ();
 sg13g2_fill_1 FILLER_66_356 ();
 sg13g2_decap_4 FILLER_66_362 ();
 sg13g2_fill_1 FILLER_66_371 ();
 sg13g2_fill_2 FILLER_66_377 ();
 sg13g2_fill_1 FILLER_66_379 ();
 sg13g2_decap_8 FILLER_66_386 ();
 sg13g2_decap_8 FILLER_66_401 ();
 sg13g2_fill_1 FILLER_66_408 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_decap_8 FILLER_67_14 ();
 sg13g2_decap_4 FILLER_67_21 ();
 sg13g2_fill_2 FILLER_67_46 ();
 sg13g2_fill_1 FILLER_67_48 ();
 sg13g2_fill_2 FILLER_67_92 ();
 sg13g2_fill_1 FILLER_67_106 ();
 sg13g2_decap_4 FILLER_67_119 ();
 sg13g2_fill_1 FILLER_67_123 ();
 sg13g2_fill_2 FILLER_67_138 ();
 sg13g2_fill_2 FILLER_67_159 ();
 sg13g2_fill_1 FILLER_67_161 ();
 sg13g2_fill_1 FILLER_67_168 ();
 sg13g2_fill_2 FILLER_67_186 ();
 sg13g2_fill_2 FILLER_67_207 ();
 sg13g2_decap_8 FILLER_67_212 ();
 sg13g2_decap_8 FILLER_67_219 ();
 sg13g2_decap_8 FILLER_67_226 ();
 sg13g2_decap_4 FILLER_67_233 ();
 sg13g2_decap_4 FILLER_67_262 ();
 sg13g2_fill_2 FILLER_67_266 ();
 sg13g2_fill_1 FILLER_67_290 ();
 sg13g2_fill_1 FILLER_67_310 ();
 sg13g2_fill_2 FILLER_67_352 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_fill_2 FILLER_67_385 ();
 sg13g2_fill_1 FILLER_67_387 ();
 sg13g2_decap_8 FILLER_67_400 ();
 sg13g2_fill_2 FILLER_67_407 ();
 sg13g2_decap_8 FILLER_68_0 ();
 sg13g2_decap_8 FILLER_68_7 ();
 sg13g2_decap_8 FILLER_68_14 ();
 sg13g2_fill_1 FILLER_68_21 ();
 sg13g2_decap_4 FILLER_68_38 ();
 sg13g2_fill_1 FILLER_68_55 ();
 sg13g2_decap_8 FILLER_68_94 ();
 sg13g2_decap_4 FILLER_68_101 ();
 sg13g2_fill_1 FILLER_68_105 ();
 sg13g2_decap_4 FILLER_68_110 ();
 sg13g2_fill_2 FILLER_68_114 ();
 sg13g2_decap_4 FILLER_68_129 ();
 sg13g2_fill_1 FILLER_68_146 ();
 sg13g2_fill_2 FILLER_68_176 ();
 sg13g2_fill_1 FILLER_68_178 ();
 sg13g2_fill_2 FILLER_68_188 ();
 sg13g2_decap_8 FILLER_68_206 ();
 sg13g2_decap_8 FILLER_68_213 ();
 sg13g2_decap_8 FILLER_68_220 ();
 sg13g2_decap_8 FILLER_68_227 ();
 sg13g2_fill_2 FILLER_68_246 ();
 sg13g2_decap_8 FILLER_68_264 ();
 sg13g2_decap_4 FILLER_68_271 ();
 sg13g2_fill_2 FILLER_68_275 ();
 sg13g2_decap_4 FILLER_68_306 ();
 sg13g2_fill_1 FILLER_68_322 ();
 sg13g2_fill_2 FILLER_68_329 ();
 sg13g2_fill_2 FILLER_68_350 ();
 sg13g2_decap_8 FILLER_68_370 ();
 sg13g2_decap_8 FILLER_68_377 ();
 sg13g2_decap_8 FILLER_68_384 ();
 sg13g2_decap_8 FILLER_68_400 ();
 sg13g2_fill_2 FILLER_68_407 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_fill_1 FILLER_69_21 ();
 sg13g2_fill_1 FILLER_69_48 ();
 sg13g2_decap_4 FILLER_69_70 ();
 sg13g2_fill_1 FILLER_69_74 ();
 sg13g2_fill_1 FILLER_69_87 ();
 sg13g2_decap_8 FILLER_69_94 ();
 sg13g2_decap_4 FILLER_69_105 ();
 sg13g2_fill_2 FILLER_69_109 ();
 sg13g2_fill_1 FILLER_69_115 ();
 sg13g2_fill_2 FILLER_69_120 ();
 sg13g2_decap_8 FILLER_69_126 ();
 sg13g2_fill_2 FILLER_69_133 ();
 sg13g2_fill_1 FILLER_69_135 ();
 sg13g2_fill_2 FILLER_69_144 ();
 sg13g2_fill_1 FILLER_69_146 ();
 sg13g2_fill_2 FILLER_69_164 ();
 sg13g2_fill_1 FILLER_69_185 ();
 sg13g2_fill_2 FILLER_69_204 ();
 sg13g2_fill_1 FILLER_69_206 ();
 sg13g2_fill_2 FILLER_69_260 ();
 sg13g2_fill_2 FILLER_69_268 ();
 sg13g2_decap_8 FILLER_69_298 ();
 sg13g2_fill_1 FILLER_69_310 ();
 sg13g2_decap_4 FILLER_69_346 ();
 sg13g2_fill_2 FILLER_69_356 ();
 sg13g2_fill_1 FILLER_69_358 ();
 sg13g2_decap_4 FILLER_69_365 ();
 sg13g2_fill_1 FILLER_69_375 ();
 sg13g2_decap_8 FILLER_69_401 ();
 sg13g2_fill_1 FILLER_69_408 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_fill_2 FILLER_70_28 ();
 sg13g2_fill_1 FILLER_70_30 ();
 sg13g2_decap_4 FILLER_70_36 ();
 sg13g2_fill_1 FILLER_70_40 ();
 sg13g2_decap_8 FILLER_70_50 ();
 sg13g2_decap_8 FILLER_70_57 ();
 sg13g2_decap_4 FILLER_70_64 ();
 sg13g2_fill_1 FILLER_70_68 ();
 sg13g2_fill_1 FILLER_70_75 ();
 sg13g2_decap_8 FILLER_70_80 ();
 sg13g2_fill_2 FILLER_70_103 ();
 sg13g2_decap_8 FILLER_70_132 ();
 sg13g2_decap_8 FILLER_70_139 ();
 sg13g2_decap_8 FILLER_70_151 ();
 sg13g2_fill_2 FILLER_70_212 ();
 sg13g2_fill_1 FILLER_70_214 ();
 sg13g2_fill_2 FILLER_70_222 ();
 sg13g2_fill_2 FILLER_70_232 ();
 sg13g2_decap_8 FILLER_70_257 ();
 sg13g2_decap_8 FILLER_70_264 ();
 sg13g2_decap_8 FILLER_70_271 ();
 sg13g2_fill_2 FILLER_70_278 ();
 sg13g2_fill_1 FILLER_70_280 ();
 sg13g2_fill_1 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_317 ();
 sg13g2_decap_8 FILLER_70_324 ();
 sg13g2_fill_2 FILLER_70_342 ();
 sg13g2_fill_2 FILLER_70_354 ();
 sg13g2_decap_8 FILLER_70_397 ();
 sg13g2_decap_4 FILLER_70_404 ();
 sg13g2_fill_1 FILLER_70_408 ();
 sg13g2_decap_8 FILLER_71_0 ();
 sg13g2_decap_8 FILLER_71_7 ();
 sg13g2_decap_8 FILLER_71_14 ();
 sg13g2_decap_8 FILLER_71_21 ();
 sg13g2_decap_8 FILLER_71_28 ();
 sg13g2_fill_1 FILLER_71_35 ();
 sg13g2_decap_8 FILLER_71_40 ();
 sg13g2_decap_8 FILLER_71_47 ();
 sg13g2_fill_1 FILLER_71_67 ();
 sg13g2_decap_4 FILLER_71_80 ();
 sg13g2_decap_8 FILLER_71_125 ();
 sg13g2_decap_8 FILLER_71_132 ();
 sg13g2_decap_8 FILLER_71_139 ();
 sg13g2_decap_8 FILLER_71_146 ();
 sg13g2_fill_1 FILLER_71_153 ();
 sg13g2_fill_1 FILLER_71_181 ();
 sg13g2_fill_1 FILLER_71_208 ();
 sg13g2_fill_1 FILLER_71_229 ();
 sg13g2_decap_8 FILLER_71_246 ();
 sg13g2_decap_4 FILLER_71_253 ();
 sg13g2_fill_2 FILLER_71_257 ();
 sg13g2_decap_4 FILLER_71_267 ();
 sg13g2_fill_2 FILLER_71_271 ();
 sg13g2_fill_1 FILLER_71_304 ();
 sg13g2_decap_8 FILLER_71_348 ();
 sg13g2_fill_2 FILLER_71_355 ();
 sg13g2_decap_8 FILLER_71_367 ();
 sg13g2_fill_2 FILLER_71_374 ();
 sg13g2_decap_8 FILLER_71_388 ();
 sg13g2_decap_8 FILLER_71_395 ();
 sg13g2_decap_8 FILLER_71_402 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_fill_2 FILLER_72_21 ();
 sg13g2_fill_1 FILLER_72_23 ();
 sg13g2_decap_4 FILLER_72_47 ();
 sg13g2_fill_2 FILLER_72_51 ();
 sg13g2_decap_4 FILLER_72_66 ();
 sg13g2_fill_2 FILLER_72_70 ();
 sg13g2_fill_2 FILLER_72_80 ();
 sg13g2_fill_1 FILLER_72_82 ();
 sg13g2_fill_1 FILLER_72_91 ();
 sg13g2_decap_4 FILLER_72_118 ();
 sg13g2_decap_8 FILLER_72_134 ();
 sg13g2_decap_8 FILLER_72_141 ();
 sg13g2_decap_4 FILLER_72_148 ();
 sg13g2_fill_1 FILLER_72_152 ();
 sg13g2_decap_4 FILLER_72_158 ();
 sg13g2_fill_2 FILLER_72_169 ();
 sg13g2_decap_8 FILLER_72_212 ();
 sg13g2_decap_8 FILLER_72_219 ();
 sg13g2_decap_8 FILLER_72_226 ();
 sg13g2_decap_8 FILLER_72_233 ();
 sg13g2_decap_8 FILLER_72_240 ();
 sg13g2_fill_1 FILLER_72_247 ();
 sg13g2_fill_2 FILLER_72_265 ();
 sg13g2_fill_2 FILLER_72_287 ();
 sg13g2_fill_1 FILLER_72_289 ();
 sg13g2_fill_2 FILLER_72_306 ();
 sg13g2_fill_1 FILLER_72_308 ();
 sg13g2_fill_2 FILLER_72_316 ();
 sg13g2_decap_4 FILLER_72_348 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_fill_2 FILLER_72_406 ();
 sg13g2_fill_1 FILLER_72_408 ();
 sg13g2_decap_8 FILLER_73_0 ();
 sg13g2_decap_8 FILLER_73_7 ();
 sg13g2_fill_2 FILLER_73_14 ();
 sg13g2_fill_1 FILLER_73_16 ();
 sg13g2_decap_8 FILLER_73_59 ();
 sg13g2_decap_4 FILLER_73_78 ();
 sg13g2_fill_2 FILLER_73_98 ();
 sg13g2_fill_1 FILLER_73_100 ();
 sg13g2_fill_2 FILLER_73_106 ();
 sg13g2_fill_1 FILLER_73_112 ();
 sg13g2_fill_1 FILLER_73_143 ();
 sg13g2_fill_2 FILLER_73_178 ();
 sg13g2_decap_8 FILLER_73_202 ();
 sg13g2_decap_8 FILLER_73_209 ();
 sg13g2_fill_2 FILLER_73_216 ();
 sg13g2_fill_1 FILLER_73_218 ();
 sg13g2_decap_4 FILLER_73_247 ();
 sg13g2_fill_1 FILLER_73_256 ();
 sg13g2_decap_8 FILLER_73_281 ();
 sg13g2_decap_8 FILLER_73_288 ();
 sg13g2_decap_8 FILLER_73_295 ();
 sg13g2_fill_2 FILLER_73_302 ();
 sg13g2_fill_2 FILLER_73_334 ();
 sg13g2_decap_4 FILLER_73_349 ();
 sg13g2_fill_2 FILLER_73_373 ();
 sg13g2_fill_1 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_4 FILLER_73_403 ();
 sg13g2_fill_2 FILLER_73_407 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_fill_2 FILLER_74_43 ();
 sg13g2_decap_4 FILLER_74_79 ();
 sg13g2_fill_2 FILLER_74_83 ();
 sg13g2_fill_2 FILLER_74_97 ();
 sg13g2_fill_1 FILLER_74_99 ();
 sg13g2_fill_2 FILLER_74_108 ();
 sg13g2_fill_1 FILLER_74_144 ();
 sg13g2_fill_1 FILLER_74_161 ();
 sg13g2_decap_8 FILLER_74_173 ();
 sg13g2_fill_1 FILLER_74_180 ();
 sg13g2_decap_8 FILLER_74_184 ();
 sg13g2_decap_8 FILLER_74_191 ();
 sg13g2_decap_8 FILLER_74_198 ();
 sg13g2_fill_1 FILLER_74_205 ();
 sg13g2_fill_2 FILLER_74_247 ();
 sg13g2_fill_1 FILLER_74_263 ();
 sg13g2_fill_2 FILLER_74_274 ();
 sg13g2_fill_2 FILLER_74_281 ();
 sg13g2_decap_4 FILLER_74_293 ();
 sg13g2_decap_8 FILLER_74_301 ();
 sg13g2_fill_1 FILLER_74_308 ();
 sg13g2_decap_8 FILLER_74_318 ();
 sg13g2_fill_2 FILLER_74_325 ();
 sg13g2_decap_8 FILLER_74_332 ();
 sg13g2_fill_2 FILLER_74_350 ();
 sg13g2_fill_1 FILLER_74_352 ();
 sg13g2_fill_2 FILLER_74_359 ();
 sg13g2_fill_2 FILLER_74_374 ();
 sg13g2_decap_8 FILLER_74_389 ();
 sg13g2_decap_8 FILLER_74_396 ();
 sg13g2_decap_4 FILLER_74_403 ();
 sg13g2_fill_2 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_fill_2 FILLER_75_28 ();
 sg13g2_fill_1 FILLER_75_30 ();
 sg13g2_fill_2 FILLER_75_36 ();
 sg13g2_fill_2 FILLER_75_47 ();
 sg13g2_fill_1 FILLER_75_49 ();
 sg13g2_decap_8 FILLER_75_71 ();
 sg13g2_decap_8 FILLER_75_78 ();
 sg13g2_fill_2 FILLER_75_98 ();
 sg13g2_fill_1 FILLER_75_100 ();
 sg13g2_fill_2 FILLER_75_105 ();
 sg13g2_fill_2 FILLER_75_111 ();
 sg13g2_fill_2 FILLER_75_120 ();
 sg13g2_decap_8 FILLER_75_130 ();
 sg13g2_decap_8 FILLER_75_166 ();
 sg13g2_decap_8 FILLER_75_173 ();
 sg13g2_decap_8 FILLER_75_180 ();
 sg13g2_decap_8 FILLER_75_187 ();
 sg13g2_fill_2 FILLER_75_194 ();
 sg13g2_fill_1 FILLER_75_239 ();
 sg13g2_fill_2 FILLER_75_268 ();
 sg13g2_fill_1 FILLER_75_280 ();
 sg13g2_fill_2 FILLER_75_304 ();
 sg13g2_fill_1 FILLER_75_311 ();
 sg13g2_decap_8 FILLER_75_316 ();
 sg13g2_decap_8 FILLER_75_323 ();
 sg13g2_decap_4 FILLER_75_330 ();
 sg13g2_fill_1 FILLER_75_334 ();
 sg13g2_decap_8 FILLER_75_338 ();
 sg13g2_decap_8 FILLER_75_345 ();
 sg13g2_fill_1 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_372 ();
 sg13g2_decap_8 FILLER_75_379 ();
 sg13g2_decap_8 FILLER_75_386 ();
 sg13g2_decap_8 FILLER_75_393 ();
 sg13g2_decap_8 FILLER_75_400 ();
 sg13g2_fill_2 FILLER_75_407 ();
 sg13g2_decap_8 FILLER_76_0 ();
 sg13g2_decap_8 FILLER_76_7 ();
 sg13g2_decap_8 FILLER_76_14 ();
 sg13g2_decap_8 FILLER_76_21 ();
 sg13g2_decap_8 FILLER_76_28 ();
 sg13g2_decap_8 FILLER_76_35 ();
 sg13g2_decap_8 FILLER_76_42 ();
 sg13g2_decap_8 FILLER_76_49 ();
 sg13g2_fill_2 FILLER_76_56 ();
 sg13g2_decap_4 FILLER_76_71 ();
 sg13g2_decap_4 FILLER_76_80 ();
 sg13g2_fill_2 FILLER_76_89 ();
 sg13g2_fill_2 FILLER_76_96 ();
 sg13g2_fill_2 FILLER_76_126 ();
 sg13g2_fill_1 FILLER_76_128 ();
 sg13g2_decap_4 FILLER_76_133 ();
 sg13g2_fill_1 FILLER_76_137 ();
 sg13g2_decap_8 FILLER_76_162 ();
 sg13g2_decap_8 FILLER_76_169 ();
 sg13g2_fill_2 FILLER_76_176 ();
 sg13g2_fill_2 FILLER_76_218 ();
 sg13g2_fill_1 FILLER_76_301 ();
 sg13g2_fill_2 FILLER_76_342 ();
 sg13g2_decap_8 FILLER_76_352 ();
 sg13g2_decap_8 FILLER_76_359 ();
 sg13g2_decap_8 FILLER_76_366 ();
 sg13g2_decap_8 FILLER_76_373 ();
 sg13g2_decap_8 FILLER_76_380 ();
 sg13g2_decap_8 FILLER_76_387 ();
 sg13g2_decap_8 FILLER_76_394 ();
 sg13g2_decap_8 FILLER_76_401 ();
 sg13g2_fill_1 FILLER_76_408 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_4 FILLER_77_49 ();
 sg13g2_fill_2 FILLER_77_98 ();
 sg13g2_fill_2 FILLER_77_108 ();
 sg13g2_fill_1 FILLER_77_110 ();
 sg13g2_fill_2 FILLER_77_128 ();
 sg13g2_decap_4 FILLER_77_143 ();
 sg13g2_decap_8 FILLER_77_152 ();
 sg13g2_decap_8 FILLER_77_159 ();
 sg13g2_decap_8 FILLER_77_166 ();
 sg13g2_decap_8 FILLER_77_173 ();
 sg13g2_fill_2 FILLER_77_180 ();
 sg13g2_fill_1 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_187 ();
 sg13g2_decap_8 FILLER_77_194 ();
 sg13g2_decap_4 FILLER_77_209 ();
 sg13g2_fill_1 FILLER_77_213 ();
 sg13g2_fill_2 FILLER_77_246 ();
 sg13g2_fill_1 FILLER_77_281 ();
 sg13g2_fill_1 FILLER_77_319 ();
 sg13g2_decap_8 FILLER_77_375 ();
 sg13g2_decap_8 FILLER_77_382 ();
 sg13g2_decap_8 FILLER_77_389 ();
 sg13g2_decap_8 FILLER_77_396 ();
 sg13g2_decap_4 FILLER_77_403 ();
 sg13g2_fill_2 FILLER_77_407 ();
 sg13g2_decap_8 FILLER_78_0 ();
 sg13g2_decap_8 FILLER_78_7 ();
 sg13g2_decap_8 FILLER_78_14 ();
 sg13g2_decap_8 FILLER_78_21 ();
 sg13g2_decap_8 FILLER_78_28 ();
 sg13g2_decap_8 FILLER_78_35 ();
 sg13g2_decap_8 FILLER_78_42 ();
 sg13g2_decap_8 FILLER_78_49 ();
 sg13g2_fill_2 FILLER_78_56 ();
 sg13g2_fill_1 FILLER_78_58 ();
 sg13g2_fill_2 FILLER_78_87 ();
 sg13g2_fill_1 FILLER_78_89 ();
 sg13g2_decap_8 FILLER_78_155 ();
 sg13g2_decap_8 FILLER_78_162 ();
 sg13g2_decap_8 FILLER_78_169 ();
 sg13g2_decap_8 FILLER_78_176 ();
 sg13g2_decap_8 FILLER_78_183 ();
 sg13g2_decap_8 FILLER_78_190 ();
 sg13g2_decap_8 FILLER_78_197 ();
 sg13g2_decap_8 FILLER_78_204 ();
 sg13g2_decap_4 FILLER_78_211 ();
 sg13g2_fill_1 FILLER_78_215 ();
 sg13g2_fill_1 FILLER_78_247 ();
 sg13g2_fill_2 FILLER_78_278 ();
 sg13g2_fill_1 FILLER_78_280 ();
 sg13g2_fill_1 FILLER_78_297 ();
 sg13g2_decap_8 FILLER_78_373 ();
 sg13g2_decap_8 FILLER_78_380 ();
 sg13g2_decap_8 FILLER_78_387 ();
 sg13g2_decap_8 FILLER_78_394 ();
 sg13g2_decap_8 FILLER_78_401 ();
 sg13g2_fill_1 FILLER_78_408 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_decap_8 FILLER_79_56 ();
 sg13g2_decap_4 FILLER_79_63 ();
 sg13g2_fill_2 FILLER_79_67 ();
 sg13g2_decap_4 FILLER_79_82 ();
 sg13g2_fill_1 FILLER_79_86 ();
 sg13g2_decap_4 FILLER_79_92 ();
 sg13g2_fill_2 FILLER_79_113 ();
 sg13g2_fill_1 FILLER_79_123 ();
 sg13g2_fill_2 FILLER_79_129 ();
 sg13g2_decap_8 FILLER_79_144 ();
 sg13g2_decap_8 FILLER_79_151 ();
 sg13g2_decap_8 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_172 ();
 sg13g2_decap_8 FILLER_79_179 ();
 sg13g2_decap_8 FILLER_79_186 ();
 sg13g2_decap_8 FILLER_79_193 ();
 sg13g2_decap_8 FILLER_79_200 ();
 sg13g2_decap_8 FILLER_79_207 ();
 sg13g2_decap_4 FILLER_79_214 ();
 sg13g2_fill_1 FILLER_79_218 ();
 sg13g2_fill_2 FILLER_79_269 ();
 sg13g2_fill_1 FILLER_79_271 ();
 sg13g2_fill_1 FILLER_79_286 ();
 sg13g2_fill_1 FILLER_79_320 ();
 sg13g2_fill_2 FILLER_79_343 ();
 sg13g2_decap_8 FILLER_79_373 ();
 sg13g2_decap_8 FILLER_79_380 ();
 sg13g2_decap_8 FILLER_79_387 ();
 sg13g2_decap_8 FILLER_79_394 ();
 sg13g2_decap_8 FILLER_79_401 ();
 sg13g2_fill_1 FILLER_79_408 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_4 FILLER_80_60 ();
 sg13g2_decap_4 FILLER_80_68 ();
 sg13g2_decap_4 FILLER_80_76 ();
 sg13g2_decap_4 FILLER_80_84 ();
 sg13g2_decap_4 FILLER_80_92 ();
 sg13g2_decap_4 FILLER_80_100 ();
 sg13g2_decap_4 FILLER_80_108 ();
 sg13g2_decap_4 FILLER_80_116 ();
 sg13g2_decap_4 FILLER_80_124 ();
 sg13g2_fill_2 FILLER_80_132 ();
 sg13g2_fill_2 FILLER_80_142 ();
 sg13g2_decap_4 FILLER_80_148 ();
 sg13g2_decap_4 FILLER_80_156 ();
 sg13g2_decap_4 FILLER_80_164 ();
 sg13g2_decap_4 FILLER_80_172 ();
 sg13g2_decap_8 FILLER_80_180 ();
 sg13g2_decap_8 FILLER_80_187 ();
 sg13g2_decap_8 FILLER_80_194 ();
 sg13g2_decap_8 FILLER_80_201 ();
 sg13g2_decap_8 FILLER_80_208 ();
 sg13g2_decap_8 FILLER_80_215 ();
 sg13g2_decap_8 FILLER_80_222 ();
 sg13g2_decap_4 FILLER_80_229 ();
 sg13g2_fill_2 FILLER_80_233 ();
 sg13g2_fill_2 FILLER_80_244 ();
 sg13g2_fill_1 FILLER_80_246 ();
 sg13g2_fill_2 FILLER_80_311 ();
 sg13g2_fill_2 FILLER_80_333 ();
 sg13g2_fill_2 FILLER_80_366 ();
 sg13g2_decap_8 FILLER_80_373 ();
 sg13g2_decap_8 FILLER_80_380 ();
 sg13g2_decap_8 FILLER_80_387 ();
 sg13g2_decap_8 FILLER_80_394 ();
 sg13g2_decap_8 FILLER_80_401 ();
 sg13g2_fill_1 FILLER_80_408 ();
 assign uio_oe[0] = net13;
 assign uio_oe[1] = net14;
 assign uio_oe[2] = net15;
 assign uio_oe[3] = net16;
 assign uio_oe[4] = net17;
 assign uio_oe[5] = net18;
 assign uio_oe[6] = net19;
 assign uio_oe[7] = net20;
 assign uio_out[0] = net21;
 assign uio_out[1] = net22;
 assign uio_out[2] = net23;
 assign uio_out[3] = net24;
 assign uio_out[4] = net25;
 assign uio_out[5] = net26;
 assign uio_out[6] = net27;
 assign uio_out[7] = net28;
endmodule
